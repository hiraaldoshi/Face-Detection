module HAAR_Comparison (



);

endmodule 