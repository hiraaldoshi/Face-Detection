module Left (

input int stage_num,
input int feature_num,
output int value

);

string name;
assign name = {"LEFT_", $sformatf("%d", stage_num), "_", $sformatf("%d", feature_num)};

always_comb
    begin

        case (name)

            "LEFT_0_0": value  <= 0.03379419073462489737;
            "LEFT_0_1": value  <= 0.15141320228576660156;
            "LEFT_0_2": value  <= 0.09004928171634669909;
            "LEFT_1_0": value  <= 0.06930858641862870650;
            "LEFT_1_1": value  <= 0.17958030104637148772;
            "LEFT_1_2": value  <= 0.16936729848384859953;
            "LEFT_1_3": value  <= 0.58663320541381835938;
            "LEFT_1_4": value  <= 0.14131669700145718660;
            "LEFT_1_5": value  <= 0.36756721138954162598;
            "LEFT_1_6": value  <= 0.61613857746124267578;
            "LEFT_1_7": value  <= 0.28362309932708740234;
            "LEFT_1_8": value  <= 0.22235809266567230225;
            "LEFT_1_9": value  <= 0.24064640700817110930;
            "LEFT_1_10": value  <= 0.55596548318862915039;
            "LEFT_1_11": value  <= 0.85027372837066650391;
            "LEFT_1_12": value  <= 0.59936738014221191406;
            "LEFT_1_13": value  <= 0.43418860435485839844;
            "LEFT_1_14": value  <= 0.30278879404067987613;
            "LEFT_1_15": value  <= 0.17984339594841000642;
            "LEFT_2_0": value  <= 0.66442251205444335938;
            "LEFT_2_1": value  <= 0.63253521919250488281;
            "LEFT_2_2": value  <= 0.12402880191802979903;
            "LEFT_2_3": value  <= 0.14321430027484891023;
            "LEFT_2_4": value  <= 0.16574330627918240633;
            "LEFT_2_5": value  <= 0.26955071091651922055;
            "LEFT_2_6": value  <= 0.18935389816761019621;
            "LEFT_2_7": value  <= 0.23093290627002718840;
            "LEFT_2_8": value  <= 0.27596020698547357730;
            "LEFT_2_9": value  <= 0.17325380444526669588;
            "LEFT_2_10": value  <= 0.13394099473953249846;
            "LEFT_2_11": value  <= 0.36287039518356317691;
            "LEFT_2_12": value  <= 0.09121105074882510100;
            "LEFT_2_13": value  <= 0.37151429057121282407;
            "LEFT_2_14": value  <= 0.59533137083053588867;
            "LEFT_2_15": value  <= 0.18440659344196319580;
            "LEFT_2_16": value  <= 0.35942441225051879883;
            "LEFT_2_17": value  <= 0.59943532943725585938;
            "LEFT_2_18": value  <= 0.41726520657539367676;
            "LEFT_2_19": value  <= 0.45097151398658752441;
            "LEFT_2_20": value  <= 0.54382127523422241211;
            "LEFT_3_0": value  <= 0.14152669906616210938;
            "LEFT_3_1": value  <= 0.61910742521286010742;
            "LEFT_3_2": value  <= 0.14873969554901120271;
            "LEFT_3_3": value  <= 0.27469098567962652035;
            "LEFT_3_4": value  <= 0.58708512783050537109;
            "LEFT_3_5": value  <= 0.58809447288513183594;
            "LEFT_3_6": value  <= 0.23733270168304440584;
            "LEFT_3_7": value  <= 0.12206549942493440108;
            "LEFT_3_8": value  <= 0.26312309503555297852;
            "LEFT_3_9": value  <= 0.36386200785636901855;
            "LEFT_3_10": value  <= 0.43035310506820678711;
            "LEFT_3_11": value  <= 0.21226030588150018863;
            "LEFT_3_12": value  <= 0.56318491697311401367;
            "LEFT_3_13": value  <= 0.57971078157424926758;
            "LEFT_3_14": value  <= 0.27052420377731317691;
            "LEFT_3_15": value  <= 0.54356247186660766602;
            "LEFT_3_16": value  <= 0.53194248676300048828;
            "LEFT_3_17": value  <= 0.54189807176589965820;
            "LEFT_3_18": value  <= 0.36953729391098022461;
            "LEFT_3_19": value  <= 0.35650369524955749512;
            "LEFT_3_20": value  <= 0.19139820337295529451;
            "LEFT_3_21": value  <= 0.38355550169944757632;
            "LEFT_3_22": value  <= 0.43128961324691772461;
            "LEFT_3_23": value  <= 0.39848309755325317383;
            "LEFT_3_24": value  <= 0.23667329549789428711;
            "LEFT_3_25": value  <= 0.58175009489059448242;
            "LEFT_3_26": value  <= 0.55405938625335693359;
            "LEFT_3_27": value  <= 0.17752550542354580965;
            "LEFT_3_28": value  <= 0.30241701006889337711;
            "LEFT_3_29": value  <= 0.44149309396743768863;
            "LEFT_3_30": value  <= 0.27913948893547058105;
            "LEFT_3_31": value  <= 0.52631992101669311523;
            "LEFT_3_32": value  <= 0.43193790316581731625;
            "LEFT_3_33": value  <= 0.30820429325103759766;
            "LEFT_3_34": value  <= 0.55219221115112304688;
            "LEFT_3_35": value  <= 0.54013228416442871094;
            "LEFT_3_36": value  <= 0.51786178350448608398;
            "LEFT_3_37": value  <= 0.52902942895889282227;
            "LEFT_3_38": value  <= 0.74719941616058349609;
            "LEFT_4_0": value  <= 0.20640860497951510344;
            "LEFT_4_1": value  <= 0.58519971370697021484;
            "LEFT_4_2": value  <= 0.09401842951774599944;
            "LEFT_4_3": value  <= 0.17819879949092870541;
            "LEFT_4_4": value  <= 0.16383990645408630371;
            "LEFT_4_5": value  <= 0.20854400098323819246;
            "LEFT_4_6": value  <= 0.57027608156204223633;
            "LEFT_4_7": value  <= 0.51169431209564208984;
            "LEFT_4_8": value  <= 0.71313798427581787109;
            "LEFT_4_9": value  <= 0.25671818852424621582;
            "LEFT_4_10": value  <= 0.17006659507751470395;
            "LEFT_4_11": value  <= 0.54105567932128906250;
            "LEFT_4_12": value  <= 0.37324368953704828433;
            "LEFT_4_13": value  <= 0.26264819502830510922;
            "LEFT_4_14": value  <= 0.20037539303302770444;
            "LEFT_4_15": value  <= 0.55919027328491210938;
            "LEFT_4_16": value  <= 0.27304071187973022461;
            "LEFT_4_17": value  <= 0.14059090614318850432;
            "LEFT_4_18": value  <= 0.17950350046157839690;
            "LEFT_4_19": value  <= 0.57367831468582153320;
            "LEFT_4_20": value  <= 0.23706759512424468994;
            "LEFT_4_21": value  <= 0.56081998348236083984;
            "LEFT_4_22": value  <= 0.16401059925556180086;
            "LEFT_4_23": value  <= 0.52276492118835449219;
            "LEFT_4_24": value  <= 0.70161938667297363281;
            "LEFT_4_25": value  <= 0.27673470973968511410;
            "LEFT_4_26": value  <= 0.43422400951385498047;
            "LEFT_4_27": value  <= 0.57264858484268188477;
            "LEFT_4_28": value  <= 0.21068480610847470369;
            "LEFT_4_29": value  <= 0.75937908887863159180;
            "LEFT_4_30": value  <= 0.12524759769439700041;
            "LEFT_4_31": value  <= 0.33153840899467468262;
            "LEFT_4_32": value  <= 0.55060499906539916992;
            "LEFT_5_0": value  <= 0.17626909911632540617;
            "LEFT_5_1": value  <= 0.61181068420410156250;
            "LEFT_5_2": value  <= 0.09904426336288449373;
            "LEFT_5_3": value  <= 0.55798798799514770508;
            "LEFT_5_4": value  <= 0.22314579784870150481;
            "LEFT_5_5": value  <= 0.26539939641952520200;
            "LEFT_5_6": value  <= 0.58038270473480224609;
            "LEFT_5_7": value  <= 0.18303519487380978670;
            "LEFT_5_8": value  <= 0.33635589480400091000;
            "LEFT_5_9": value  <= 0.22866420447826391049;
            "LEFT_5_10": value  <= 0.56259131431579589844;
            "LEFT_5_11": value  <= 0.39069938659667968750;
            "LEFT_5_12": value  <= 0.52484822273254394531;
            "LEFT_5_13": value  <= 0.41943109035491937808;
            "LEFT_5_14": value  <= 0.18825499713420870695;
            "LEFT_5_15": value  <= 0.13399730622768399324;
            "LEFT_5_16": value  <= 0.37620881199836730957;
            "LEFT_5_17": value  <= 0.26631429791450500488;
            "LEFT_5_18": value  <= 0.53635787963867187500;
            "LEFT_5_19": value  <= 0.53582328557968139648;
            "LEFT_5_20": value  <= 0.24096719920635220613;
            "LEFT_5_21": value  <= 0.54258567094802856445;
            "LEFT_5_22": value  <= 0.41584059596061712094;
            "LEFT_5_23": value  <= 0.28112530708312988281;
            "LEFT_5_24": value  <= 0.52600282430648803711;
            "LEFT_5_25": value  <= 0.56735092401504516602;
            "LEFT_5_26": value  <= 0.53435921669006347656;
            "LEFT_5_27": value  <= 0.60108900070190429688;
            "LEFT_5_28": value  <= 0.81991511583328247070;
            "LEFT_5_29": value  <= 0.22002810239791870117;
            "LEFT_5_30": value  <= 0.44130811095237731934;
            "LEFT_5_31": value  <= 0.54788607358932495117;
            "LEFT_5_32": value  <= 0.63578677177429199219;
            "LEFT_5_33": value  <= 0.34936860203742980957;
            "LEFT_5_34": value  <= 0.11196149885654449463;
            "LEFT_5_35": value  <= 0.23871029913425451108;
            "LEFT_5_36": value  <= 0.75869178771972656250;
            "LEFT_5_37": value  <= 0.25654768943786621094;
            "LEFT_5_38": value  <= 0.67343479394912719727;
            "LEFT_5_39": value  <= 0.54883527755737304688;
            "LEFT_5_40": value  <= 0.61043310165405273438;
            "LEFT_5_41": value  <= 0.53108531236648559570;
            "LEFT_5_42": value  <= 0.17291119694709780608;
            "LEFT_5_43": value  <= 0.65977597236633300781;
            "LEFT_6_0": value  <= 0.61034351587295532227;
            "LEFT_6_1": value  <= 0.26323631405830377750;
            "LEFT_6_2": value  <= 0.58728742599487304688;
            "LEFT_6_3": value  <= 0.15678019821643829346;
            "LEFT_6_4": value  <= 0.19131539762020111084;
            "LEFT_6_5": value  <= 0.29149138927459722348;
            "LEFT_6_6": value  <= 0.19434769451618200131;
            "LEFT_6_7": value  <= 0.31346169114112848453;
            "LEFT_6_8": value  <= 0.25364819169044500180;
            "LEFT_6_9": value  <= 0.57677221298217773438;
            "LEFT_6_10": value  <= 0.28431910276412958316;
            "LEFT_6_11": value  <= 0.40524271130561828613;
            "LEFT_6_12": value  <= 0.57837551832199096680;
            "LEFT_6_13": value  <= 0.55413120985031127930;
            "LEFT_6_14": value  <= 0.40326559543609619141;
            "LEFT_6_15": value  <= 0.35359779000282287598;
            "LEFT_6_16": value  <= 0.30374449491500848941;
            "LEFT_6_17": value  <= 0.71810871362686157227;
            "LEFT_6_18": value  <= 0.56219518184661865234;
            "LEFT_6_19": value  <= 0.46153879165649408511;
            "LEFT_6_20": value  <= 0.53438371419906616211;
            "LEFT_6_21": value  <= 0.16862459480762478914;
            "LEFT_6_22": value  <= 0.37920561432838439941;
            "LEFT_6_23": value  <= 0.15128670632839200105;
            "LEFT_6_24": value  <= 0.20818220078945159912;
            "LEFT_6_25": value  <= 0.40982469916343688965;
            "LEFT_6_26": value  <= 0.56932741403579711914;
            "LEFT_6_27": value  <= 0.53267508745193481445;
            "LEFT_6_28": value  <= 0.15513050556182861328;
            "LEFT_6_29": value  <= 0.55005669593811035156;
            "LEFT_6_30": value  <= 0.42386838793754577637;
            "LEFT_6_31": value  <= 0.21500380337238308992;
            "LEFT_6_32": value  <= 0.66757112741470336914;
            "LEFT_6_33": value  <= 0.22672890126705169678;
            "LEFT_6_34": value  <= 0.43086910247802728824;
            "LEFT_6_35": value  <= 0.58366149663925170898;
            "LEFT_6_36": value  <= 0.70169448852539062500;
            "LEFT_6_37": value  <= 0.28953450918197631836;
            "LEFT_6_38": value  <= 0.29755708575248718262;
            "LEFT_6_39": value  <= 0.48888179659843450375;
            "LEFT_6_40": value  <= 0.14814929664134979248;
            "LEFT_6_41": value  <= 0.47863098978996282407;
            "LEFT_6_42": value  <= 0.73742228746414184570;
            "LEFT_6_43": value  <= 0.34891548752784729004;
            "LEFT_6_44": value  <= 0.23796869814395910092;
            "LEFT_6_45": value  <= 0.19646880030632019043;
            "LEFT_6_46": value  <= 0.55905228853225708008;
            "LEFT_6_47": value  <= 0.06340465694665910201;
            "LEFT_6_48": value  <= 0.73234677314758300781;
            "LEFT_6_49": value  <= 0.41148349642753601074;
            "LEFT_7_0": value  <= 0.26635450124740600586;
            "LEFT_7_1": value  <= 0.61438488960266113281;
            "LEFT_7_2": value  <= 0.57663410902023315430;
            "LEFT_7_3": value  <= 0.56820458173751831055;
            "LEFT_7_4": value  <= 0.16406759619712829590;
            "LEFT_7_5": value  <= 0.61231541633605957031;
            "LEFT_7_6": value  <= 0.57078588008880615234;
            "LEFT_7_7": value  <= 0.40896728634834289551;
            "LEFT_7_8": value  <= 0.57124507427215576172;
            "LEFT_7_9": value  <= 0.52625042200088500977;
            "LEFT_7_10": value  <= 0.68538308143615722656;
            "LEFT_7_11": value  <= 0.32662820816040039062;
            "LEFT_7_12": value  <= 0.54684108495712280273;
            "LEFT_7_13": value  <= 0.55706679821014404297;
            "LEFT_7_14": value  <= 0.37005689740180969238;
            "LEFT_7_15": value  <= 0.21400700509548190031;
            "LEFT_7_16": value  <= 0.55267721414566040039;
            "LEFT_7_17": value  <= 0.39580118656158447266;
            "LEFT_7_18": value  <= 0.52413737773895263672;
            "LEFT_7_19": value  <= 0.33854091167449951172;
            "LEFT_7_20": value  <= 0.54853779077529907227;
            "LEFT_7_21": value  <= 0.33752760291099548340;
            "LEFT_7_22": value  <= 0.56317430734634399414;
            "LEFT_7_23": value  <= 0.06373503804206849532;
            "LEFT_7_24": value  <= 0.51369631290435791016;
            "LEFT_7_25": value  <= 0.38793200254440307617;
            "LEFT_7_26": value  <= 0.52500867843627929688;
            "LEFT_7_27": value  <= 0.66720288991928100586;
            "LEFT_7_28": value  <= 0.71633791923522949219;
            "LEFT_7_29": value  <= 0.30213609337806701660;
            "LEFT_7_30": value  <= 0.18200090527534490414;
            "LEFT_7_31": value  <= 0.33891880512237548828;
            "LEFT_7_32": value  <= 0.40853491425514221191;
            "LEFT_7_33": value  <= 0.33783990144729608707;
            "LEFT_7_34": value  <= 0.42046359181404108218;
            "LEFT_7_35": value  <= 0.25952160358428960629;
            "LEFT_7_36": value  <= 0.61651438474655151367;
            "LEFT_7_37": value  <= 0.16280280053615570068;
            "LEFT_7_38": value  <= 0.31996509432792658023;
            "LEFT_7_39": value  <= 0.41039940714836120605;
            "LEFT_7_40": value  <= 0.10349129885435100207;
            "LEFT_7_41": value  <= 0.84938651323318481445;
            "LEFT_7_42": value  <= 0.31301578879356378726;
            "LEFT_7_43": value  <= 0.48563209176063537598;
            "LEFT_7_44": value  <= 0.83946740627288818359;
            "LEFT_7_45": value  <= 0.18816959857940671053;
            "LEFT_7_46": value  <= 0.52712291479110717773;
            "LEFT_7_47": value  <= 0.42353048920631408691;
            "LEFT_7_48": value  <= 0.69343960285186767578;
            "LEFT_7_49": value  <= 0.59009212255477905273;
            "LEFT_7_50": value  <= 0.64663827419281005859;
            "LEFT_8_0": value  <= 0.61423242092132568359;
            "LEFT_8_1": value  <= 0.57049518823623657227;
            "LEFT_8_2": value  <= 0.21122519671916958894;
            "LEFT_8_3": value  <= 0.29504820704460138492;
            "LEFT_8_4": value  <= 0.29909908771514892578;
            "LEFT_8_5": value  <= 0.28130298852920532227;
            "LEFT_8_6": value  <= 0.35353690385818481445;
            "LEFT_8_7": value  <= 0.55965322256088256836;
            "LEFT_8_8": value  <= 0.59780317544937133789;
            "LEFT_8_9": value  <= 0.27552521228790277652;
            "LEFT_8_10": value  <= 0.43056419491767877750;
            "LEFT_8_11": value  <= 0.24952429533004760742;
            "LEFT_8_12": value  <= 0.54785531759262084961;
            "LEFT_8_13": value  <= 0.39386010169982910156;
            "LEFT_8_14": value  <= 0.44076061248779302426;
            "LEFT_8_15": value  <= 0.54452431201934814453;
            "LEFT_8_16": value  <= 0.25447669625282287598;
            "LEFT_8_17": value  <= 0.27188581228256231137;
            "LEFT_8_18": value  <= 0.31782880425453191586;
            "LEFT_8_19": value  <= 0.42842191457748407535;
            "LEFT_8_20": value  <= 0.59028607606887817383;
            "LEFT_8_21": value  <= 0.38164898753166198730;
            "LEFT_8_22": value  <= 0.17477439343929290771;
            "LEFT_8_23": value  <= 0.36017221212387090512;
            "LEFT_8_24": value  <= 0.54018580913543701172;
            "LEFT_8_25": value  <= 0.32207700610160827637;
            "LEFT_8_26": value  <= 0.43015280365943908691;
            "LEFT_8_27": value  <= 0.35645830631256097965;
            "LEFT_8_28": value  <= 0.34907829761505132504;
            "LEFT_8_29": value  <= 0.17762720584869390317;
            "LEFT_8_30": value  <= 0.61496877670288085938;
            "LEFT_8_31": value  <= 0.54130148887634277344;
            "LEFT_8_32": value  <= 0.64494907855987548828;
            "LEFT_8_33": value  <= 0.54001551866531372070;
            "LEFT_8_34": value  <= 0.27745240926742548160;
            "LEFT_8_35": value  <= 0.56767392158508300781;
            "LEFT_8_36": value  <= 0.77492219209671020508;
            "LEFT_8_37": value  <= 0.53387218713760375977;
            "LEFT_8_38": value  <= 0.56119632720947265625;
            "LEFT_8_39": value  <= 0.29152289032936101743;
            "LEFT_8_40": value  <= 0.55364328622817993164;
            "LEFT_8_41": value  <= 0.37543910741806030273;
            "LEFT_8_42": value  <= 0.70196992158889770508;
            "LEFT_8_43": value  <= 0.23103649914264678955;
            "LEFT_8_44": value  <= 0.58648687601089477539;
            "LEFT_8_45": value  <= 0.37324070930480962582;
            "LEFT_8_46": value  <= 0.53120911121368408203;
            "LEFT_8_47": value  <= 0.47100159525871282407;
            "LEFT_8_48": value  <= 0.51678192615509033203;
            "LEFT_8_49": value  <= 0.53976088762283325195;
            "LEFT_8_50": value  <= 0.70864880084991455078;
            "LEFT_8_51": value  <= 0.52064812183380126953;
            "LEFT_8_52": value  <= 0.35070759057998657227;
            "LEFT_8_53": value  <= 0.58595228195190429688;
            "LEFT_8_54": value  <= 0.67432671785354614258;
            "LEFT_8_55": value  <= 0.52827161550521850586;
            "LEFT_9_0": value  <= 0.59147310256958007812;
            "LEFT_9_1": value  <= 0.23125819861888891049;
            "LEFT_9_2": value  <= 0.16565300524234768953;
            "LEFT_9_3": value  <= 0.54234498739242553711;
            "LEFT_9_4": value  <= 0.34179040789604192563;
            "LEFT_9_5": value  <= 0.37195819616317749023;
            "LEFT_9_6": value  <= 0.25774860382080078125;
            "LEFT_9_7": value  <= 0.29507490992546081543;
            "LEFT_9_8": value  <= 0.75693589448928833008;
            "LEFT_9_9": value  <= 0.55837088823318481445;
            "LEFT_9_10": value  <= 0.56273132562637329102;
            "LEFT_9_11": value  <= 0.27711850404739379883;
            "LEFT_9_12": value  <= 0.55806517601013183594;
            "LEFT_9_13": value  <= 0.33302500844001770020;
            "LEFT_9_14": value  <= 0.29905349016189580746;
            "LEFT_9_15": value  <= 0.14638589322566988860;
            "LEFT_9_16": value  <= 0.37469539046287542172;
            "LEFT_9_17": value  <= 0.27547478675842290707;
            "LEFT_9_18": value  <= 0.37445840239524841309;
            "LEFT_9_19": value  <= 0.75138592720031738281;
            "LEFT_9_20": value  <= 0.54048967361450195312;
            "LEFT_9_21": value  <= 0.61697798967361450195;
            "LEFT_9_22": value  <= 0.20484960079193120785;
            "LEFT_9_23": value  <= 0.52529847621917724609;
            "LEFT_9_24": value  <= 0.52677828073501586914;
            "LEFT_9_25": value  <= 0.69545578956604003906;
            "LEFT_9_26": value  <= 0.42918878793716430664;
            "LEFT_9_27": value  <= 0.29305368661880487613;
            "LEFT_9_28": value  <= 0.44953250885009771176;
            "LEFT_9_29": value  <= 0.31491199135780328922;
            "LEFT_9_30": value  <= 0.51218920946121215820;
            "LEFT_9_31": value  <= 0.51759117841720581055;
            "LEFT_9_32": value  <= 0.51371401548385620117;
            "LEFT_9_33": value  <= 0.55743098258972167969;
            "LEFT_9_34": value  <= 0.55489408969879150391;
            "LEFT_9_35": value  <= 0.33874198794364929199;
            "LEFT_9_36": value  <= 0.53580617904663085938;
            "LEFT_9_37": value  <= 0.61252027750015258789;
            "LEFT_9_38": value  <= 0.23581659793853759766;
            "LEFT_9_39": value  <= 0.73231112957000732422;
            "LEFT_9_40": value  <= 0.54194551706314086914;
            "LEFT_9_41": value  <= 0.28216940164566040039;
            "LEFT_9_42": value  <= 0.91299301385879516602;
            "LEFT_9_43": value  <= 0.60226702690124511719;
            "LEFT_9_44": value  <= 0.56132131814956665039;
            "LEFT_9_45": value  <= 0.22616119682788848877;
            "LEFT_9_46": value  <= 0.40756919980049127750;
            "LEFT_9_47": value  <= 0.28272539377212518863;
            "LEFT_9_48": value  <= 0.50747412443161010742;
            "LEFT_9_49": value  <= 0.61690068244934082031;
            "LEFT_9_50": value  <= 0.45244330167770391293;
            "LEFT_9_51": value  <= 0.52404087781906127930;
            "LEFT_9_52": value  <= 0.52093791961669921875;
            "LEFT_9_53": value  <= 0.54507029056549072266;
            "LEFT_9_54": value  <= 0.69990468025207519531;
            "LEFT_9_55": value  <= 0.26536649465560907535;
            "LEFT_9_56": value  <= 0.44805660843849182129;
            "LEFT_9_57": value  <= 0.42313501238822942563;
            "LEFT_9_58": value  <= 0.53417021036148071289;
            "LEFT_9_59": value  <= 0.51186597347259521484;
            "LEFT_9_60": value  <= 0.35321870446205139160;
            "LEFT_9_61": value  <= 0.28423538804054260254;
            "LEFT_9_62": value  <= 0.68836402893066406250;
            "LEFT_9_63": value  <= 0.17098939418792730160;
            "LEFT_9_64": value  <= 0.52908462285995483398;
            "LEFT_9_65": value  <= 0.64988541603088378906;
            "LEFT_9_66": value  <= 0.32604381442070007324;
            "LEFT_9_67": value  <= 0.75289410352706909180;
            "LEFT_9_68": value  <= 0.53351658582687377930;
            "LEFT_9_69": value  <= 0.45803940296173101254;
            "LEFT_9_70": value  <= 0.25923201441764831543;
            "LEFT_10_0": value  <= 0.32588860392570501157;
            "LEFT_10_1": value  <= 0.58388811349868774414;
            "LEFT_10_2": value  <= 0.57080817222595214844;
            "LEFT_10_3": value  <= 0.25010511279106140137;
            "LEFT_10_4": value  <= 0.23853680491447448730;
            "LEFT_10_5": value  <= 0.39550709724426269531;
            "LEFT_10_6": value  <= 0.56397080421447753906;
            "LEFT_10_7": value  <= 0.21865129470825200864;
            "LEFT_10_8": value  <= 0.23507060110569000244;
            "LEFT_10_9": value  <= 0.38041129708290100098;
            "LEFT_10_10": value  <= 0.25101679563522338867;
            "LEFT_10_11": value  <= 0.59928238391876220703;
            "LEFT_10_12": value  <= 0.56813961267471313477;
            "LEFT_10_13": value  <= 0.14913170039653780852;
            "LEFT_10_14": value  <= 0.36924299597740167789;
            "LEFT_10_15": value  <= 0.67585092782974243164;
            "LEFT_10_16": value  <= 0.53680229187011718750;
            "LEFT_10_17": value  <= 0.16493770480155950375;
            "LEFT_10_18": value  <= 0.19639259576797490903;
            "LEFT_10_19": value  <= 0.46711719036102300473;
            "LEFT_10_20": value  <= 0.11554169654846190018;
            "LEFT_10_21": value  <= 0.51496601104736328125;
            "LEFT_10_22": value  <= 0.36054810881614690610;
            "LEFT_10_23": value  <= 0.48862120509147638492;
            "LEFT_10_24": value  <= 0.53568130731582641602;
            "LEFT_10_25": value  <= 0.18486219644546508789;
            "LEFT_10_26": value  <= 0.38405799865722661801;
            "LEFT_10_27": value  <= 0.42885640263557428531;
            "LEFT_10_28": value  <= 0.29136741161346441098;
            "LEFT_10_29": value  <= 0.75547999143600463867;
            "LEFT_10_30": value  <= 0.28382799029350280762;
            "LEFT_10_31": value  <= 0.48709350824356079102;
            "LEFT_10_32": value  <= 0.70997077226638793945;
            "LEFT_10_33": value  <= 0.40308868885040277652;
            "LEFT_10_34": value  <= 0.45020240545272832700;
            "LEFT_10_35": value  <= 0.54428607225418090820;
            "LEFT_10_36": value  <= 0.42004638910293579102;
            "LEFT_10_37": value  <= 0.37925618886947631836;
            "LEFT_10_38": value  <= 0.72531038522720336914;
            "LEFT_10_39": value  <= 0.46933019161224370785;
            "LEFT_10_40": value  <= 0.51492130756378173828;
            "LEFT_10_41": value  <= 0.53997439146041870117;
            "LEFT_10_42": value  <= 0.24084959924221038818;
            "LEFT_10_43": value  <= 0.65735882520675659180;
            "LEFT_10_44": value  <= 0.41928219795227050781;
            "LEFT_10_45": value  <= 0.55402982234954833984;
            "LEFT_10_46": value  <= 0.17109179496765139494;
            "LEFT_10_47": value  <= 0.19042180478572851010;
            "LEFT_10_48": value  <= 0.44475069642066961118;
            "LEFT_10_49": value  <= 0.24907270073890688811;
            "LEFT_10_50": value  <= 0.53812432289123535156;
            "LEFT_10_51": value  <= 0.55302321910858154297;
            "LEFT_10_52": value  <= 0.41326990723609918765;
            "LEFT_10_53": value  <= 0.09878723323345180163;
            "LEFT_10_54": value  <= 0.09112749248743060027;
            "LEFT_10_55": value  <= 0.47266489267349237613;
            "LEFT_10_56": value  <= 0.21574570238590240479;
            "LEFT_10_57": value  <= 0.54107707738876342773;
            "LEFT_10_58": value  <= 0.77878749370574951172;
            "LEFT_10_59": value  <= 0.54789870977401733398;
            "LEFT_10_60": value  <= 0.53305608034133911133;
            "LEFT_10_61": value  <= 0.69235211610794067383;
            "LEFT_10_62": value  <= 0.50559002161026000977;
            "LEFT_10_63": value  <= 0.37837418913841247559;
            "LEFT_10_64": value  <= 0.30816510319709777832;
            "LEFT_10_65": value  <= 0.66339588165283203125;
            "LEFT_10_66": value  <= 0.65968447923660278320;
            "LEFT_10_67": value  <= 0.52318328619003295898;
            "LEFT_10_68": value  <= 0.52042502164840698242;
            "LEFT_10_69": value  <= 0.72388780117034912109;
            "LEFT_10_70": value  <= 0.31050220131874078922;
            "LEFT_10_71": value  <= 0.31389680504798889160;
            "LEFT_10_72": value  <= 0.45365801453590387515;
            "LEFT_10_73": value  <= 0.18044540286064150725;
            "LEFT_10_74": value  <= 0.72557020187377929688;
            "LEFT_10_75": value  <= 0.44129210710525512695;
            "LEFT_10_76": value  <= 0.35000529885292047672;
            "LEFT_10_77": value  <= 0.49121949076652532407;
            "LEFT_10_78": value  <= 0.35702759027481079102;
            "LEFT_10_79": value  <= 0.43537721037864690610;
            "LEFT_11_0": value  <= 0.61625832319259643555;
            "LEFT_11_1": value  <= 0.58182948827743530273;
            "LEFT_11_2": value  <= 0.25520521402359008789;
            "LEFT_11_3": value  <= 0.36850899457931518555;
            "LEFT_11_4": value  <= 0.23323920369148248843;
            "LEFT_11_5": value  <= 0.32574570178985601254;
            "LEFT_11_6": value  <= 0.37447169423103332520;
            "LEFT_11_7": value  <= 0.34203711152076721191;
            "LEFT_11_8": value  <= 0.28044199943542480469;
            "LEFT_11_9": value  <= 0.25790509581565862485;
            "LEFT_11_10": value  <= 0.41751560568809509277;
            "LEFT_11_11": value  <= 0.58651697635650634766;
            "LEFT_11_12": value  <= 0.52111411094665527344;
            "LEFT_11_13": value  <= 0.27534329891204828433;
            "LEFT_11_14": value  <= 0.57229787111282348633;
            "LEFT_11_15": value  <= 0.44661080837249761410;
            "LEFT_11_16": value  <= 0.28132531046867370605;
            "LEFT_11_17": value  <= 0.43997099995613098145;
            "LEFT_11_18": value  <= 0.29811179637908941098;
            "LEFT_11_19": value  <= 0.77052152156829833984;
            "LEFT_11_20": value  <= 0.37188440561294561215;
            "LEFT_11_21": value  <= 0.36151960492134088687;
            "LEFT_11_22": value  <= 0.53647047281265258789;
            "LEFT_11_23": value  <= 0.69276517629623413086;
            "LEFT_11_24": value  <= 0.77121537923812866211;
            "LEFT_11_25": value  <= 0.33749839663505548648;
            "LEFT_11_26": value  <= 0.53251898288726806641;
            "LEFT_11_27": value  <= 0.68376529216766357422;
            "LEFT_11_28": value  <= 0.35720878839492797852;
            "LEFT_11_29": value  <= 0.55414271354675292969;
            "LEFT_11_30": value  <= 0.50708442926406860352;
            "LEFT_11_31": value  <= 0.52695602178573608398;
            "LEFT_11_32": value  <= 0.71455889940261840820;
            "LEFT_11_33": value  <= 0.53986120223999023438;
            "LEFT_11_34": value  <= 0.24391929805278780852;
            "LEFT_11_35": value  <= 0.38868919014930730649;
            "LEFT_11_36": value  <= 0.33894580602645868472;
            "LEFT_11_37": value  <= 0.46014139056205749512;
            "LEFT_11_38": value  <= 0.57698792219161987305;
            "LEFT_11_39": value  <= 0.48787090182304382324;
            "LEFT_11_40": value  <= 0.52635532617568969727;
            "LEFT_11_41": value  <= 0.14988289773464200105;
            "LEFT_11_42": value  <= 0.02489331923425200030;
            "LEFT_11_43": value  <= 0.54646229743957519531;
            "LEFT_11_44": value  <= 0.42710569500923162289;
            "LEFT_11_45": value  <= 0.68741792440414428711;
            "LEFT_11_46": value  <= 0.33706760406494140625;
            "LEFT_11_47": value  <= 0.46267929673194890805;
            "LEFT_11_48": value  <= 0.53461229801177978516;
            "LEFT_11_49": value  <= 0.46438300609588617496;
            "LEFT_11_50": value  <= 0.51963961124420166016;
            "LEFT_11_51": value  <= 0.48381629586219787598;
            "LEFT_11_52": value  <= 0.89203029870986938477;
            "LEFT_11_53": value  <= 0.20339429378509518709;
            "LEFT_11_54": value  <= 0.45716339349746698550;
            "LEFT_11_55": value  <= 0.52711081504821777344;
            "LEFT_11_56": value  <= 0.41383129358291631528;
            "LEFT_11_57": value  <= 0.52251511812210083008;
            "LEFT_11_58": value  <= 0.52367687225341796875;
            "LEFT_11_59": value  <= 0.45310598611831670590;
            "LEFT_11_60": value  <= 0.51308518648147583008;
            "LEFT_11_61": value  <= 0.77865952253341674805;
            "LEFT_11_62": value  <= 0.42885988950729370117;
            "LEFT_11_63": value  <= 0.35239779949188232422;
            "LEFT_11_64": value  <= 0.68410861492156982422;
            "LEFT_11_65": value  <= 0.35655200481414800473;
            "LEFT_11_66": value  <= 0.33687931299209600278;
            "LEFT_11_67": value  <= 0.34221610426902770996;
            "LEFT_11_68": value  <= 0.65336120128631591797;
            "LEFT_11_69": value  <= 0.53075802326202392578;
            "LEFT_11_70": value  <= 0.68574589490890502930;
            "LEFT_11_71": value  <= 0.40378510951995849609;
            "LEFT_11_72": value  <= 0.53997987508773803711;
            "LEFT_11_73": value  <= 0.46654370427131647281;
            "LEFT_11_74": value  <= 0.59147810935974121094;
            "LEFT_11_75": value  <= 0.36420381069183349609;
            "LEFT_11_76": value  <= 0.26642319560050958804;
            "LEFT_11_77": value  <= 0.67795312404632568359;
            "LEFT_11_78": value  <= 0.56139647960662841797;
            "LEFT_11_79": value  <= 0.59644782543182373047;
            "LEFT_11_80": value  <= 0.29761150479316711426;
            "LEFT_11_81": value  <= 0.51878392696380615234;
            "LEFT_11_82": value  <= 0.18660229444503778629;
            "LEFT_11_83": value  <= 0.52121251821517944336;
            "LEFT_11_84": value  <= 0.45899370312690740414;
            "LEFT_11_85": value  <= 0.30799409747123718262;
            "LEFT_11_86": value  <= 0.21010440587997439299;
            "LEFT_11_87": value  <= 0.57653552293777465820;
            "LEFT_11_88": value  <= 0.50651001930236816406;
            "LEFT_11_89": value  <= 0.49669149518013000488;
            "LEFT_11_90": value  <= 0.21949790418148040771;
            "LEFT_11_91": value  <= 0.47784018516540527344;
            "LEFT_11_92": value  <= 0.19363629817962649260;
            "LEFT_11_93": value  <= 0.59990632534027099609;
            "LEFT_11_94": value  <= 0.33383339643478388004;
            "LEFT_11_95": value  <= 0.66170698404312133789;
            "LEFT_11_96": value  <= 0.44887441396713262387;
            "LEFT_11_97": value  <= 0.54093921184539794922;
            "LEFT_11_98": value  <= 0.68191200494766235352;
            "LEFT_11_99": value  <= 0.46307921409606928043;
            "LEFT_11_100": value  <= 0.51653790473937988281;
            "LEFT_11_101": value  <= 0.25363931059837341309;
            "LEFT_11_102": value  <= 0.39851561188697820493;
            "LEFT_12_0": value  <= 0.28910180926322942563;
            "LEFT_12_1": value  <= 0.62117892503738403320;
            "LEFT_12_2": value  <= 0.22544120252132421323;
            "LEFT_12_3": value  <= 0.37117108702659612485;
            "LEFT_12_4": value  <= 0.56517201662063598633;
            "LEFT_12_5": value  <= 0.30691260099411010742;
            "LEFT_12_6": value  <= 0.57628279924392700195;
            "LEFT_12_7": value  <= 0.26442441344261169434;
            "LEFT_12_8": value  <= 0.50511389970779418945;
            "LEFT_12_9": value  <= 0.58269691467285156250;
            "LEFT_12_10": value  <= 0.31138521432876592465;
            "LEFT_12_11": value  <= 0.32779461145401000977;
            "LEFT_12_12": value  <= 0.73817098140716552734;
            "LEFT_12_13": value  <= 0.52566307783126831055;
            "LEFT_12_14": value  <= 0.55112308263778686523;
            "LEFT_12_15": value  <= 0.54256367683410644531;
            "LEFT_12_16": value  <= 0.53801918029785156250;
            "LEFT_12_17": value  <= 0.30358019471168518066;
            "LEFT_12_18": value  <= 0.39909970760345458984;
            "LEFT_12_19": value  <= 0.55628067255020141602;
            "LEFT_12_20": value  <= 0.46096539497375488281;
            "LEFT_12_21": value  <= 0.23161660134792330656;
            "LEFT_12_22": value  <= 0.23307719826698300447;
            "LEFT_12_23": value  <= 0.46574440598487848453;
            "LEFT_12_24": value  <= 0.51543921232223510742;
            "LEFT_12_25": value  <= 0.62197732925415039062;
            "LEFT_12_26": value  <= 0.18373550474643710051;
            "LEFT_12_27": value  <= 0.51459872722625732422;
            "LEFT_12_28": value  <= 0.53436601161956787109;
            "LEFT_12_29": value  <= 0.62150079011917114258;
            "LEFT_12_30": value  <= 0.42992618680000310727;
            "LEFT_12_31": value  <= 0.52603340148925781250;
            "LEFT_12_32": value  <= 0.35065388679504400082;
            "LEFT_12_33": value  <= 0.48096409440040588379;
            "LEFT_12_34": value  <= 0.11393620073795319991;
            "LEFT_12_35": value  <= 0.63520950078964233398;
            "LEFT_12_36": value  <= 0.51311182975769042969;
            "LEFT_12_37": value  <= 0.54213947057723999023;
            "LEFT_12_38": value  <= 0.18949599564075469971;
            "LEFT_12_39": value  <= 0.64543670415878295898;
            "LEFT_12_40": value  <= 0.62150311470031738281;
            "LEFT_12_41": value  <= 0.37126109004020690918;
            "LEFT_12_42": value  <= 0.50236439704895019531;
            "LEFT_12_43": value  <= 0.32402679324150091000;
            "LEFT_12_44": value  <= 0.41655078530311578922;
            "LEFT_12_45": value  <= 0.38540428876876831055;
            "LEFT_12_46": value  <= 0.22044940292835241147;
            "LEFT_12_47": value  <= 0.56070661544799804688;
            "LEFT_12_48": value  <= 0.46216571331024169922;
            "LEFT_12_49": value  <= 0.52695941925048828125;
            "LEFT_12_50": value  <= 0.63592231273651123047;
            "LEFT_12_51": value  <= 0.52747678756713867188;
            "LEFT_12_52": value  <= 0.20385199785232541170;
            "LEFT_12_53": value  <= 0.45874550938606262207;
            "LEFT_12_54": value  <= 0.50712740421295166016;
            "LEFT_12_55": value  <= 0.48121041059494018555;
            "LEFT_12_56": value  <= 0.46258139610290527344;
            "LEFT_12_57": value  <= 0.53862917423248291016;
            "LEFT_12_58": value  <= 0.02594250068068500170;
            "LEFT_12_59": value  <= 0.52028447389602661133;
            "LEFT_12_60": value  <= 0.72824811935424804688;
            "LEFT_12_61": value  <= 0.55623567104339599609;
            "LEFT_12_62": value  <= 0.68033927679061889648;
            "LEFT_12_63": value  <= 0.25616711378097528629;
            "LEFT_12_64": value  <= 0.51896202564239501953;
            "LEFT_12_65": value  <= 0.12950749695301058684;
            "LEFT_12_66": value  <= 0.57350981235504150391;
            "LEFT_12_67": value  <= 0.52898782491683959961;
            "LEFT_12_68": value  <= 0.65756398439407348633;
            "LEFT_12_69": value  <= 0.36280471086502080746;
            "LEFT_12_70": value  <= 0.12842659652233121004;
            "LEFT_12_71": value  <= 0.62922400236129760742;
            "LEFT_12_72": value  <= 0.14877319335937500000;
            "LEFT_12_73": value  <= 0.42561021447181701660;
            "LEFT_12_74": value  <= 0.40041440725326538086;
            "LEFT_12_75": value  <= 0.60091161727905273438;
            "LEFT_12_76": value  <= 0.35149338841438287906;
            "LEFT_12_77": value  <= 0.46422758698463439941;
            "LEFT_12_78": value  <= 0.50255292654037475586;
            "LEFT_12_79": value  <= 0.58845919370651245117;
            "LEFT_12_80": value  <= 0.43722391128540039062;
            "LEFT_12_81": value  <= 0.43275511264801030942;
            "LEFT_12_82": value  <= 0.19131340086460110750;
            "LEFT_12_83": value  <= 0.53081780672073364258;
            "LEFT_12_84": value  <= 0.63653957843780517578;
            "LEFT_12_85": value  <= 0.51898342370986938477;
            "LEFT_12_86": value  <= 0.51050621271133422852;
            "LEFT_12_87": value  <= 0.46969148516654968262;
            "LEFT_12_88": value  <= 0.50536459684371948242;
            "LEFT_12_89": value  <= 0.65089809894561767578;
            "LEFT_12_90": value  <= 0.62418168783187866211;
            "LEFT_12_91": value  <= 0.34327811002731317691;
            "LEFT_12_92": value  <= 0.18780590593814849854;
            "LEFT_12_93": value  <= 0.38052770495414728336;
            "LEFT_12_94": value  <= 0.68437147140502929688;
            "LEFT_12_95": value  <= 0.55029052495956420898;
            "LEFT_12_96": value  <= 0.33688580989837652035;
            "LEFT_12_97": value  <= 0.64876401424407958984;
            "LEFT_12_98": value  <= 0.40345790982246398926;
            "LEFT_12_99": value  <= 0.63868737220764160156;
            "LEFT_12_100": value  <= 0.29864218831062322446;
            "LEFT_12_101": value  <= 0.50221997499465942383;
            "LEFT_12_102": value  <= 0.64924520254135131836;
            "LEFT_12_103": value  <= 0.51505708694458007812;
            "LEFT_12_104": value  <= 0.45736691355705261230;
            "LEFT_12_105": value  <= 0.38655120134353637695;
            "LEFT_12_106": value  <= 0.51285791397094726562;
            "LEFT_12_107": value  <= 0.40515819191932678223;
            "LEFT_12_108": value  <= 0.52959501743316650391;
            "LEFT_12_109": value  <= 0.47894069552421569824;
            "LEFT_12_110": value  <= 0.53844892978668212891;
            "LEFT_13_0": value  <= 0.39485278725624078922;
            "LEFT_13_1": value  <= 0.33703160285949712582;
            "LEFT_13_2": value  <= 0.35005760192871088199;
            "LEFT_13_3": value  <= 0.32675281167030328922;
            "LEFT_13_4": value  <= 0.30445998907089227847;
            "LEFT_13_5": value  <= 0.36500120162963872739;
            "LEFT_13_6": value  <= 0.33135411143302917480;
            "LEFT_13_7": value  <= 0.26979428529739379883;
            "LEFT_13_8": value  <= 0.52693581581115722656;
            "LEFT_13_9": value  <= 0.29096031188964838199;
            "LEFT_13_10": value  <= 0.58925771713256835938;
            "LEFT_13_11": value  <= 0.35235640406608581543;
            "LEFT_13_12": value  <= 0.54230177402496337891;
            "LEFT_13_13": value  <= 0.51939457654953002930;
            "LEFT_13_14": value  <= 0.31577691435813898257;
            "LEFT_13_15": value  <= 0.44512999057769780942;
            "LEFT_13_16": value  <= 0.30317419767379760742;
            "LEFT_13_17": value  <= 0.47814530134201049805;
            "LEFT_13_18": value  <= 0.31863081455230707340;
            "LEFT_13_19": value  <= 0.64135968685150146484;
            "LEFT_13_20": value  <= 0.15074980258941650391;
            "LEFT_13_21": value  <= 0.43161588907241821289;
            "LEFT_13_22": value  <= 0.47355538606643682309;
            "LEFT_13_23": value  <= 0.35531890392303472348;
            "LEFT_13_24": value  <= 0.45000949501991271973;
            "LEFT_13_25": value  <= 0.56292420625686645508;
            "LEFT_13_26": value  <= 0.53815472126007080078;
            "LEFT_13_27": value  <= 0.52559971809387207031;
            "LEFT_13_28": value  <= 0.22728569805622100830;
            "LEFT_13_29": value  <= 0.46263080835342407227;
            "LEFT_13_30": value  <= 0.63175398111343383789;
            "LEFT_13_31": value  <= 0.54211097955703735352;
            "LEFT_13_32": value  <= 0.53584778308868408203;
            "LEFT_13_33": value  <= 0.77935767173767089844;
            "LEFT_13_34": value  <= 0.52973198890686035156;
            "LEFT_13_35": value  <= 0.46780940890312200375;
            "LEFT_13_36": value  <= 0.52767342329025268555;
            "LEFT_13_37": value  <= 0.48346799612045288086;
            "LEFT_13_38": value  <= 0.45118591189384460449;
            "LEFT_13_39": value  <= 0.53356587886810302734;
            "LEFT_13_40": value  <= 0.42507070302963262387;
            "LEFT_13_41": value  <= 0.30033200979232788086;
            "LEFT_13_42": value  <= 0.50673192739486694336;
            "LEFT_13_43": value  <= 0.47950699925422668457;
            "LEFT_13_44": value  <= 0.51331132650375366211;
            "LEFT_13_45": value  <= 0.19388419389724728670;
            "LEFT_13_46": value  <= 0.56865382194519042969;
            "LEFT_13_47": value  <= 0.42241689562797551938;
            "LEFT_13_48": value  <= 0.51137751340866088867;
            "LEFT_13_49": value  <= 0.71946620941162109375;
            "LEFT_13_50": value  <= 0.38402619957923889160;
            "LEFT_13_51": value  <= 0.59370887279510498047;
            "LEFT_13_52": value  <= 0.51385760307312011719;
            "LEFT_13_53": value  <= 0.60900372266769409180;
            "LEFT_13_54": value  <= 0.34586110711097717285;
            "LEFT_13_55": value  <= 0.56931042671203613281;
            "LEFT_13_56": value  <= 0.43505370616912841797;
            "LEFT_13_57": value  <= 0.14688730239868161287;
            "LEFT_13_58": value  <= 0.52935242652893066406;
            "LEFT_13_59": value  <= 0.46524509787559509277;
            "LEFT_13_60": value  <= 0.46535089612007141113;
            "LEFT_13_61": value  <= 0.54972952604293823242;
            "LEFT_13_62": value  <= 0.39190879464149480649;
            "LEFT_13_63": value  <= 0.16313570737838750668;
            "LEFT_13_64": value  <= 0.51458978652954101562;
            "LEFT_13_65": value  <= 0.65176361799240112305;
            "LEFT_13_66": value  <= 0.55146527290344238281;
            "LEFT_13_67": value  <= 0.31652408838272100278;
            "LEFT_13_68": value  <= 0.68533778190612792969;
            "LEFT_13_69": value  <= 0.54845881462097167969;
            "LEFT_13_70": value  <= 0.63957798480987548828;
            "LEFT_13_71": value  <= 0.27510729432106018066;
            "LEFT_13_72": value  <= 0.33256360888481140137;
            "LEFT_13_73": value  <= 0.59422808885574340820;
            "LEFT_13_74": value  <= 0.41671109199523931332;
            "LEFT_13_75": value  <= 0.54338949918746948242;
            "LEFT_13_76": value  <= 0.64071899652481079102;
            "LEFT_13_77": value  <= 0.52145552635192871094;
            "LEFT_13_78": value  <= 0.31515279412269592285;
            "LEFT_13_79": value  <= 0.48708370327949518375;
            "LEFT_13_80": value  <= 0.35697489976882940121;
            "LEFT_13_81": value  <= 0.88259208202362060547;
            "LEFT_13_82": value  <= 0.14461620151996609773;
            "LEFT_13_83": value  <= 0.53964787721633911133;
            "LEFT_13_84": value  <= 0.41704109311103820801;
            "LEFT_13_85": value  <= 0.46983671188354492188;
            "LEFT_13_86": value  <= 0.62677729129791259766;
            "LEFT_13_87": value  <= 0.30970111489295959473;
            "LEFT_13_88": value  <= 0.08112388849258420076;
            "LEFT_13_89": value  <= 0.51555037498474121094;
            "LEFT_13_90": value  <= 0.46997779607772832700;
            "LEFT_13_91": value  <= 0.39205300807952880859;
            "LEFT_13_92": value  <= 0.52606582641601562500;
            "LEFT_13_93": value  <= 0.63392949104309082031;
            "LEFT_13_94": value  <= 0.53330272436141967773;
            "LEFT_13_95": value  <= 0.17653420567512509431;
            "LEFT_13_96": value  <= 0.53241598606109619141;
            "LEFT_13_97": value  <= 0.46479299664497381039;
            "LEFT_13_98": value  <= 0.32367089390754699707;
            "LEFT_13_99": value  <= 0.47874391078948980160;
            "LEFT_13_100": value  <= 0.44093081355094909668;
            "LEFT_13_101": value  <= 0.40381139516830438785;
            "LEFT_14_0": value  <= 0.66001719236373901367;
            "LEFT_14_1": value  <= 0.57839912176132202148;
            "LEFT_14_2": value  <= 0.36222669482231140137;
            "LEFT_14_3": value  <= 0.55004191398620605469;
            "LEFT_14_4": value  <= 0.26731699705123901367;
            "LEFT_14_5": value  <= 0.38550278544425958804;
            "LEFT_14_6": value  <= 0.55032098293304443359;
            "LEFT_14_7": value  <= 0.32912218570709228516;
            "LEFT_14_8": value  <= 0.35883820056915277652;
            "LEFT_14_9": value  <= 0.42968419194221502133;
            "LEFT_14_10": value  <= 0.52821648120880126953;
            "LEFT_14_11": value  <= 0.45595678687095642090;
            "LEFT_14_12": value  <= 0.23501169681549069490;
            "LEFT_14_13": value  <= 0.53294152021408081055;
            "LEFT_14_14": value  <= 0.42730879783630371094;
            "LEFT_14_15": value  <= 0.29126119613647460938;
            "LEFT_14_16": value  <= 0.53076881170272827148;
            "LEFT_14_17": value  <= 0.47037750482559198550;
            "LEFT_14_18": value  <= 0.21415670216083529387;
            "LEFT_14_19": value  <= 0.47664138674736017398;
            "LEFT_14_20": value  <= 0.53607988357543945312;
            "LEFT_14_21": value  <= 0.57201302051544189453;
            "LEFT_14_22": value  <= 0.36931228637695312500;
            "LEFT_14_23": value  <= 0.49623748660087591000;
            "LEFT_14_24": value  <= 0.44389459490776062012;
            "LEFT_14_25": value  <= 0.52442502975463867188;
            "LEFT_14_26": value  <= 0.60602837800979614258;
            "LEFT_14_27": value  <= 0.38911709189414978027;
            "LEFT_14_28": value  <= 0.50693458318710327148;
            "LEFT_14_29": value  <= 0.58822017908096313477;
            "LEFT_14_30": value  <= 0.55336058139801025391;
            "LEFT_14_31": value  <= 0.33101469278335571289;
            "LEFT_14_32": value  <= 0.54338318109512329102;
            "LEFT_14_33": value  <= 0.56003582477569580078;
            "LEFT_14_34": value  <= 0.66854667663574218750;
            "LEFT_14_35": value  <= 0.53571212291717529297;
            "LEFT_14_36": value  <= 0.46798178553581237793;
            "LEFT_14_37": value  <= 0.39375010132789611816;
            "LEFT_14_38": value  <= 0.42423760890960687808;
            "LEFT_14_39": value  <= 0.36312100291252141782;
            "LEFT_14_40": value  <= 0.68604522943496704102;
            "LEFT_14_41": value  <= 0.39440968632698059082;
            "LEFT_14_42": value  <= 0.19626219570636749268;
            "LEFT_14_43": value  <= 0.40862590074539190121;
            "LEFT_14_44": value  <= 0.44891211390495300293;
            "LEFT_14_45": value  <= 0.53359258174896240234;
            "LEFT_14_46": value  <= 0.51113212108612060547;
            "LEFT_14_47": value  <= 0.55414897203445434570;
            "LEFT_14_48": value  <= 0.45864239335060119629;
            "LEFT_14_49": value  <= 0.53924250602722167969;
            "LEFT_14_50": value  <= 0.17037139832973480225;
            "LEFT_14_51": value  <= 0.53054618835449218750;
            "LEFT_14_52": value  <= 0.46155458688735961914;
            "LEFT_14_53": value  <= 0.48335990309715270996;
            "LEFT_14_54": value  <= 0.51876372098922729492;
            "LEFT_14_55": value  <= 0.40792569518089288882;
            "LEFT_14_56": value  <= 0.53316092491149902344;
            "LEFT_14_57": value  <= 0.56554222106933593750;
            "LEFT_14_58": value  <= 0.45343810319900512695;
            "LEFT_14_59": value  <= 0.53506332635879516602;
            "LEFT_14_60": value  <= 0.11136870086193090268;
            "LEFT_14_61": value  <= 0.56287378072738647461;
            "LEFT_14_62": value  <= 0.41658350825309747867;
            "LEFT_14_63": value  <= 0.48603910207748407535;
            "LEFT_14_64": value  <= 0.52623051404953002930;
            "LEFT_14_65": value  <= 0.53193771839141845703;
            "LEFT_14_66": value  <= 0.46182450652122497559;
            "LEFT_14_67": value  <= 0.55056709051132202148;
            "LEFT_14_68": value  <= 0.46978530287742620297;
            "LEFT_14_69": value  <= 0.38308390974998468570;
            "LEFT_14_70": value  <= 0.25663000345230102539;
            "LEFT_14_71": value  <= 0.64699661731719970703;
            "LEFT_14_72": value  <= 0.47459828853607177734;
            "LEFT_14_73": value  <= 0.53066647052764892578;
            "LEFT_14_74": value  <= 0.54131257534027099609;
            "LEFT_14_75": value  <= 0.61585122346878051758;
            "LEFT_14_76": value  <= 0.46958059072494512387;
            "LEFT_14_77": value  <= 0.28495660424232477359;
            "LEFT_14_78": value  <= 0.70569849014282226562;
            "LEFT_14_79": value  <= 0.39029321074485778809;
            "LEFT_14_80": value  <= 0.36842319369316101074;
            "LEFT_14_81": value  <= 0.38491758704185491391;
            "LEFT_14_82": value  <= 0.47297719120979309082;
            "LEFT_14_83": value  <= 0.48091810941696172543;
            "LEFT_14_84": value  <= 0.69036781787872314453;
            "LEFT_14_85": value  <= 0.53706902265548706055;
            "LEFT_14_86": value  <= 0.51398652791976928711;
            "LEFT_14_87": value  <= 0.46602371335029602051;
            "LEFT_14_88": value  <= 0.44048359990119928531;
            "LEFT_14_89": value  <= 0.54359710216522216797;
            "LEFT_14_90": value  <= 0.53705781698226928711;
            "LEFT_14_91": value  <= 0.56594127416610717773;
            "LEFT_14_92": value  <= 0.51616579294204711914;
            "LEFT_14_93": value  <= 0.48696619272232061215;
            "LEFT_14_94": value  <= 0.27274489402771001645;
            "LEFT_14_95": value  <= 0.68514388799667358398;
            "LEFT_14_96": value  <= 0.42844650149345397949;
            "LEFT_14_97": value  <= 0.42261189222335820981;
            "LEFT_14_98": value  <= 0.47446319460868841000;
            "LEFT_14_99": value  <= 0.42450588941574102231;
            "LEFT_14_100": value  <= 0.59523570537567138672;
            "LEFT_14_101": value  <= 0.41377940773963928223;
            "LEFT_14_102": value  <= 0.44841149449348449707;
            "LEFT_14_103": value  <= 0.56248587369918823242;
            "LEFT_14_104": value  <= 0.46377518773078918457;
            "LEFT_14_105": value  <= 0.45445030927658081055;
            "LEFT_14_106": value  <= 0.53347527980804443359;
            "LEFT_14_107": value  <= 0.53985852003097534180;
            "LEFT_14_108": value  <= 0.43178731203079218082;
            "LEFT_14_109": value  <= 0.17859250307083129883;
            "LEFT_14_110": value  <= 0.43424990773200988770;
            "LEFT_14_111": value  <= 0.51617169380187988281;
            "LEFT_14_112": value  <= 0.59867632389068603516;
            "LEFT_14_113": value  <= 0.41082179546356201172;
            "LEFT_14_114": value  <= 0.51738142967224121094;
            "LEFT_14_115": value  <= 0.68889832496643066406;
            "LEFT_14_116": value  <= 0.51785671710968017578;
            "LEFT_14_117": value  <= 0.16784210503101348877;
            "LEFT_14_118": value  <= 0.43682569265365600586;
            "LEFT_14_119": value  <= 0.78022962808609008789;
            "LEFT_14_120": value  <= 0.15851010382175451108;
            "LEFT_14_121": value  <= 0.51633048057556152344;
            "LEFT_14_122": value  <= 0.37283179163932800293;
            "LEFT_14_123": value  <= 0.58383792638778686523;
            "LEFT_14_124": value  <= 0.47282868623733520508;
            "LEFT_14_125": value  <= 0.53022021055221557617;
            "LEFT_14_126": value  <= 0.49983340501785278320;
            "LEFT_14_127": value  <= 0.05083335936069489913;
            "LEFT_14_128": value  <= 0.67981338500976562500;
            "LEFT_14_129": value  <= 0.60107719898223876953;
            "LEFT_14_130": value  <= 0.33933979272842407227;
            "LEFT_14_131": value  <= 0.43651369214057922363;
            "LEFT_14_132": value  <= 0.50527238845825195312;
            "LEFT_14_133": value  <= 0.57339739799499511719;
            "LEFT_14_134": value  <= 0.38922891020774841309;
            "LEFT_15_0": value  <= 0.32769501209259027652;
            "LEFT_15_1": value  <= 0.42564851045608520508;
            "LEFT_15_2": value  <= 0.37114870548248291016;
            "LEFT_15_3": value  <= 0.20411339402198788728;
            "LEFT_15_4": value  <= 0.54161262512207031250;
            "LEFT_15_5": value  <= 0.52778327465057373047;
            "LEFT_15_6": value  <= 0.53082311153411865234;
            "LEFT_15_7": value  <= 0.57738727331161499023;
            "LEFT_15_8": value  <= 0.43174389004707341977;
            "LEFT_15_9": value  <= 0.29339039325714111328;
            "LEFT_15_10": value  <= 0.54688447713851928711;
            "LEFT_15_11": value  <= 0.42815428972244262695;
            "LEFT_15_12": value  <= 0.37473011016845697574;
            "LEFT_15_13": value  <= 0.45377838611602777652;
            "LEFT_15_14": value  <= 0.29713419079780578613;
            "LEFT_15_15": value  <= 0.66990667581558227539;
            "LEFT_15_16": value  <= 0.33849540352821350098;
            "LEFT_15_17": value  <= 0.53991222381591796875;
            "LEFT_15_18": value  <= 0.44825780391693120785;
            "LEFT_15_19": value  <= 0.37112379074096679688;
            "LEFT_15_20": value  <= 0.60310882329940795898;
            "LEFT_15_21": value  <= 0.28387540578842157535;
            "LEFT_15_22": value  <= 0.52095472812652587891;
            "LEFT_15_23": value  <= 0.51199698448181152344;
            "LEFT_15_24": value  <= 0.33171200752258300781;
            "LEFT_15_25": value  <= 0.52475982904434204102;
            "LEFT_15_26": value  <= 0.57500940561294555664;
            "LEFT_15_27": value  <= 0.43424451351165771484;
            "LEFT_15_28": value  <= 0.45791471004486078433;
            "LEFT_15_29": value  <= 0.52743119001388549805;
            "LEFT_15_30": value  <= 0.71003687381744384766;
            "LEFT_15_31": value  <= 0.52792161703109741211;
            "LEFT_15_32": value  <= 0.50725251436233520508;
            "LEFT_15_33": value  <= 0.42831051349639892578;
            "LEFT_15_34": value  <= 0.55193877220153808594;
            "LEFT_15_35": value  <= 0.68670022487640380859;
            "LEFT_15_36": value  <= 0.37288740277290338687;
            "LEFT_15_37": value  <= 0.60601520538330078125;
            "LEFT_15_38": value  <= 0.50496357679367065430;
            "LEFT_15_39": value  <= 0.16312399506568908691;
            "LEFT_15_40": value  <= 0.44632780551910400391;
            "LEFT_15_41": value  <= 0.54733848571777343750;
            "LEFT_15_42": value  <= 0.11669850349426269531;
            "LEFT_15_43": value  <= 0.47692871093750000000;
            "LEFT_15_44": value  <= 0.34710898995399480649;
            "LEFT_15_45": value  <= 0.47852361202239990234;
            "LEFT_15_46": value  <= 0.58147960901260375977;
            "LEFT_15_47": value  <= 0.38780000805854797363;
            "LEFT_15_48": value  <= 0.16600510478019708804;
            "LEFT_15_49": value  <= 0.40933910012245178223;
            "LEFT_15_50": value  <= 0.62061947584152221680;
            "LEFT_15_51": value  <= 0.55677592754364013672;
            "LEFT_15_52": value  <= 0.56389278173446655273;
            "LEFT_15_53": value  <= 0.48262658715248107910;
            "LEFT_15_54": value  <= 0.50483798980712890625;
            "LEFT_15_55": value  <= 0.23695489764213559236;
            "LEFT_15_56": value  <= 0.50488287210464477539;
            "LEFT_15_57": value  <= 0.62386047840118408203;
            "LEFT_15_58": value  <= 0.33141419291496282407;
            "LEFT_15_59": value  <= 0.23800450563430788908;
            "LEFT_15_60": value  <= 0.40696358680725097656;
            "LEFT_15_61": value  <= 0.55067062377929687500;
            "LEFT_15_62": value  <= 0.55257099866867065430;
            "LEFT_15_63": value  <= 0.54554748535156250000;
            "LEFT_15_64": value  <= 0.51579958200454711914;
            "LEFT_15_65": value  <= 0.50132077932357788086;
            "LEFT_15_66": value  <= 0.55397182703018188477;
            "LEFT_15_67": value  <= 0.44250950217247009277;
            "LEFT_15_68": value  <= 0.71457821130752563477;
            "LEFT_15_69": value  <= 0.40704450011253362485;
            "LEFT_15_70": value  <= 0.78846907615661621094;
            "LEFT_15_71": value  <= 0.42961919307708740234;
            "LEFT_15_72": value  <= 0.46931621432304382324;
            "LEFT_15_73": value  <= 0.52423220872879028320;
            "LEFT_15_74": value  <= 0.50117397308349609375;
            "LEFT_15_75": value  <= 0.48285821080207830258;
            "LEFT_15_76": value  <= 0.59064859151840209961;
            "LEFT_15_77": value  <= 0.52410978078842163086;
            "LEFT_15_78": value  <= 0.30414658784866327457;
            "LEFT_15_79": value  <= 0.41281390190124511719;
            "LEFT_15_80": value  <= 0.58083951473236083984;
            "LEFT_15_81": value  <= 0.52465528249740600586;
            "LEFT_15_82": value  <= 0.46749550104141240903;
            "LEFT_15_83": value  <= 0.54094868898391723633;
            "LEFT_15_84": value  <= 0.37586399912834167480;
            "LEFT_15_85": value  <= 0.43295788764953607730;
            "LEFT_15_86": value  <= 0.52806180715560913086;
            "LEFT_15_87": value  <= 0.49021130800247192383;
            "LEFT_15_88": value  <= 0.55708801746368408203;
            "LEFT_15_89": value  <= 0.56584399938583374023;
            "LEFT_15_90": value  <= 0.60567390918731689453;
            "LEFT_15_91": value  <= 0.53904771804809570312;
            "LEFT_15_92": value  <= 0.43548288941383361816;
            "LEFT_15_93": value  <= 0.30109131336212158203;
            "LEFT_15_94": value  <= 0.53001511096954345703;
            "LEFT_15_95": value  <= 0.53280287981033325195;
            "LEFT_15_96": value  <= 0.54917281866073608398;
            "LEFT_15_97": value  <= 0.14407220482826230135;
            "LEFT_15_98": value  <= 0.77477252483367919922;
            "LEFT_15_99": value  <= 0.53554338216781616211;
            "LEFT_15_100": value  <= 0.57672351598739624023;
            "LEFT_15_101": value  <= 0.52156740427017211914;
            "LEFT_15_102": value  <= 0.49942049384117132016;
            "LEFT_15_103": value  <= 0.47422000765800481625;
            "LEFT_15_104": value  <= 0.53479540348052978516;
            "LEFT_15_105": value  <= 0.67271918058395385742;
            "LEFT_15_106": value  <= 0.31066751480102539062;
            "LEFT_15_107": value  <= 0.48863101005554199219;
            "LEFT_15_108": value  <= 0.60257941484451293945;
            "LEFT_15_109": value  <= 0.52407479286193847656;
            "LEFT_15_110": value  <= 0.50118672847747802734;
            "LEFT_15_111": value  <= 0.48667120933532720395;
            "LEFT_15_112": value  <= 0.34078910946846008301;
            "LEFT_15_113": value  <= 0.55755722522735595703;
            "LEFT_15_114": value  <= 0.64020007848739624023;
            "LEFT_15_115": value  <= 0.37664419412612920590;
            "LEFT_15_116": value  <= 0.33186489343643188477;
            "LEFT_15_117": value  <= 0.49035701155662542172;
            "LEFT_15_118": value  <= 0.15360510349273678865;
            "LEFT_15_119": value  <= 0.05882313102483750084;
            "LEFT_15_120": value  <= 0.69614887237548828125;
            "LEFT_15_121": value  <= 0.51679861545562744141;
            "LEFT_15_122": value  <= 0.42730781435966491699;
            "LEFT_15_123": value  <= 0.46389439702034002133;
            "LEFT_15_124": value  <= 0.53016489744186401367;
            "LEFT_15_125": value  <= 0.56306940317153930664;
            "LEFT_15_126": value  <= 0.43075358867645258121;
            "LEFT_15_127": value  <= 0.14448820054531100188;
            "LEFT_15_128": value  <= 0.43844321370124822446;
            "LEFT_15_129": value  <= 0.53404158353805541992;
            "LEFT_15_130": value  <= 0.52138561010360717773;
            "LEFT_15_131": value  <= 0.47694149613380432129;
            "LEFT_15_132": value  <= 0.42450091242790222168;
            "LEFT_15_133": value  <= 0.54577308893203735352;
            "LEFT_15_134": value  <= 0.57645887136459350586;
            "LEFT_15_135": value  <= 0.63728231191635131836;
            "LEFT_15_136": value  <= 0.53178739547729492188;
            "LEFT_16_0": value  <= 0.65555167198181152344;
            "LEFT_16_1": value  <= 0.37480720877647399902;
            "LEFT_16_2": value  <= 0.54254919290542602539;
            "LEFT_16_3": value  <= 0.24624420702457430754;
            "LEFT_16_4": value  <= 0.55943220853805541992;
            "LEFT_16_5": value  <= 0.39585039019584661313;
            "LEFT_16_6": value  <= 0.36989969015121459961;
            "LEFT_16_7": value  <= 0.37110909819602971860;
            "LEFT_16_8": value  <= 0.74927550554275512695;
            "LEFT_16_9": value  <= 0.56497871875762939453;
            "LEFT_16_10": value  <= 0.33810880780220031738;
            "LEFT_16_11": value  <= 0.55192911624908447266;
            "LEFT_16_12": value  <= 0.56082147359848022461;
            "LEFT_16_13": value  <= 0.35592061281204218082;
            "LEFT_16_14": value  <= 0.54147958755493164062;
            "LEFT_16_15": value  <= 0.63479030132293701172;
            "LEFT_16_16": value  <= 0.39134898781776428223;
            "LEFT_16_17": value  <= 0.25548928976058959961;
            "LEFT_16_18": value  <= 0.51746791601181030273;
            "LEFT_16_19": value  <= 0.53884482383728027344;
            "LEFT_16_20": value  <= 0.43360430002212518863;
            "LEFT_16_21": value  <= 0.52873617410659790039;
            "LEFT_16_22": value  <= 0.70194488763809204102;
            "LEFT_16_23": value  <= 0.29865521192550659180;
            "LEFT_16_24": value  <= 0.43234738707542419434;
            "LEFT_16_25": value  <= 0.52868640422821044922;
            "LEFT_16_26": value  <= 0.26584190130233770200;
            "LEFT_16_27": value  <= 0.54635268449783325195;
            "LEFT_16_28": value  <= 0.47034969925880432129;
            "LEFT_16_29": value  <= 0.20692589879035949707;
            "LEFT_16_30": value  <= 0.51826488971710205078;
            "LEFT_16_31": value  <= 0.68037772178649902344;
            "LEFT_16_32": value  <= 0.50583988428115844727;
            "LEFT_16_33": value  <= 0.29634249210357671567;
            "LEFT_16_34": value  <= 0.46554958820343017578;
            "LEFT_16_35": value  <= 0.47803479433059692383;
            "LEFT_16_36": value  <= 0.42869961261749267578;
            "LEFT_16_37": value  <= 0.52993071079254150391;
            "LEFT_16_38": value  <= 0.36746388673782348633;
            "LEFT_16_39": value  <= 0.23514920473098760434;
            "LEFT_16_40": value  <= 0.71159368753433227539;
            "LEFT_16_41": value  <= 0.44626510143280029297;
            "LEFT_16_42": value  <= 0.59456187486648559570;
            "LEFT_16_43": value  <= 0.53532499074935913086;
            "LEFT_16_44": value  <= 0.37602680921554570981;
            "LEFT_16_45": value  <= 0.63099128007888793945;
            "LEFT_16_46": value  <= 0.52301818132400512695;
            "LEFT_16_47": value  <= 0.51671397686004638672;
            "LEFT_16_48": value  <= 0.49794390797615051270;
            "LEFT_16_49": value  <= 0.71296507120132446289;
            "LEFT_16_50": value  <= 0.22881029546260830965;
            "LEFT_16_51": value  <= 0.46324339509010320493;
            "LEFT_16_52": value  <= 0.64674210548400878906;
            "LEFT_16_53": value  <= 0.14820009469985959139;
            "LEFT_16_54": value  <= 0.51354891061782836914;
            "LEFT_16_55": value  <= 0.27405610680580139160;
            "LEFT_16_56": value  <= 0.53326708078384399414;
            "LEFT_16_57": value  <= 0.53656041622161865234;
            "LEFT_16_58": value  <= 0.46537590026855468750;
            "LEFT_16_59": value  <= 0.54495012760162353516;
            "LEFT_16_60": value  <= 0.16560870409011840820;
            "LEFT_16_61": value  <= 0.51327311992645263672;
            "LEFT_16_62": value  <= 0.46179479360580438785;
            "LEFT_16_63": value  <= 0.59162509441375732422;
            "LEFT_16_64": value  <= 0.38884091377258300781;
            "LEFT_16_65": value  <= 0.41590648889541631528;
            "LEFT_16_66": value  <= 0.30890220403671270200;
            "LEFT_16_67": value  <= 0.39721998572349548340;
            "LEFT_16_68": value  <= 0.62574082612991333008;
            "LEFT_16_69": value  <= 0.20852099359035489168;
            "LEFT_16_70": value  <= 0.52224272489547729492;
            "LEFT_16_71": value  <= 0.58039271831512451172;
            "LEFT_16_72": value  <= 0.44012719392776489258;
            "LEFT_16_73": value  <= 0.53223252296447753906;
            "LEFT_16_74": value  <= 0.37418448925018310547;
            "LEFT_16_75": value  <= 0.46310418844223022461;
            "LEFT_16_76": value  <= 0.50446701049804687500;
            "LEFT_16_77": value  <= 0.72891211509704589844;
            "LEFT_16_78": value  <= 0.66671347618103027344;
            "LEFT_16_79": value  <= 0.43917590379714971371;
            "LEFT_16_80": value  <= 0.43464401364326482602;
            "LEFT_16_81": value  <= 0.44771409034728998355;
            "LEFT_16_82": value  <= 0.47402000427246088199;
            "LEFT_16_83": value  <= 0.53650617599487304688;
            "LEFT_16_84": value  <= 0.17522190511226651277;
            "LEFT_16_85": value  <= 0.72712367773056030273;
            "LEFT_16_86": value  <= 0.40039089322090148926;
            "LEFT_16_87": value  <= 0.56056129932403564453;
            "LEFT_16_88": value  <= 0.47532469034194951840;
            "LEFT_16_89": value  <= 0.53932619094848632812;
            "LEFT_16_90": value  <= 0.42408001422882080078;
            "LEFT_16_91": value  <= 0.42445999383926391602;
            "LEFT_16_92": value  <= 0.58958417177200317383;
            "LEFT_16_93": value  <= 0.26471349596977228336;
            "LEFT_16_94": value  <= 0.73476827144622802734;
            "LEFT_16_95": value  <= 0.27560499310493469238;
            "LEFT_16_96": value  <= 0.35105609893798828125;
            "LEFT_16_97": value  <= 0.56379258632659912109;
            "LEFT_16_98": value  <= 0.46145731210708618164;
            "LEFT_16_99": value  <= 0.29983788728713989258;
            "LEFT_16_100": value  <= 0.50778847932815551758;
            "LEFT_16_101": value  <= 0.48610189557075500488;
            "LEFT_16_102": value  <= 0.16733959317207339201;
            "LEFT_16_103": value  <= 0.26927569508552551270;
            "LEFT_16_104": value  <= 0.71838641166687011719;
            "LEFT_16_105": value  <= 0.52239668369293212891;
            "LEFT_16_106": value  <= 0.57193559408187866211;
            "LEFT_16_107": value  <= 0.54728418588638305664;
            "LEFT_16_108": value  <= 0.49738121032714838199;
            "LEFT_16_109": value  <= 0.47091740369796747379;
            "LEFT_16_110": value  <= 0.40896269679069519043;
            "LEFT_16_111": value  <= 0.61043697595596313477;
            "LEFT_16_112": value  <= 0.50696891546249389648;
            "LEFT_16_113": value  <= 0.48469170928001398257;
            "LEFT_16_114": value  <= 0.06052614003419880262;
            "LEFT_16_115": value  <= 0.53631097078323364258;
            "LEFT_16_116": value  <= 0.05966033041477199900;
            "LEFT_16_117": value  <= 0.47129771113395690918;
            "LEFT_16_118": value  <= 0.43635380268096918277;
            "LEFT_16_119": value  <= 0.58111858367919921875;
            "LEFT_16_120": value  <= 0.53117001056671142578;
            "LEFT_16_121": value  <= 0.37707018852233892270;
            "LEFT_16_122": value  <= 0.47661679983139038086;
            "LEFT_16_123": value  <= 0.52644628286361694336;
            "LEFT_16_124": value  <= 0.67371982336044311523;
            "LEFT_16_125": value  <= 0.56448352336883544922;
            "LEFT_16_126": value  <= 0.45260611176490778140;
            "LEFT_16_127": value  <= 0.60705822706222534180;
            "LEFT_16_128": value  <= 0.59982132911682128906;
            "LEFT_16_129": value  <= 0.42055889964103698730;
            "LEFT_16_130": value  <= 0.52064472436904907227;
            "LEFT_16_131": value  <= 0.31447041034698491879;
            "LEFT_16_132": value  <= 0.33801960945129400082;
            "LEFT_16_133": value  <= 0.58299607038497924805;
            "LEFT_16_134": value  <= 0.61631447076797485352;
            "LEFT_16_135": value  <= 0.51663571596145629883;
            "LEFT_16_136": value  <= 0.34080120921134948730;
            "LEFT_16_137": value  <= 0.61055189371109008789;
            "LEFT_16_138": value  <= 0.43272709846496582031;
            "LEFT_16_139": value  <= 0.48556530475616460629;
            "LEFT_17_0": value  <= 0.33325248956680297852;
            "LEFT_17_1": value  <= 0.34906411170959472656;
            "LEFT_17_2": value  <= 0.55425661802291870117;
            "LEFT_17_3": value  <= 0.36125791072845458984;
            "LEFT_17_4": value  <= 0.35301390290260320493;
            "LEFT_17_5": value  <= 0.39167788624763488770;
            "LEFT_17_6": value  <= 0.46674820780754089355;
            "LEFT_17_7": value  <= 0.30736848711967468262;
            "LEFT_17_8": value  <= 0.56221181154251098633;
            "LEFT_17_9": value  <= 0.52676612138748168945;
            "LEFT_17_10": value  <= 0.66683208942413330078;
            "LEFT_17_11": value  <= 0.55214381217956542969;
            "LEFT_17_12": value  <= 0.36286780238151550293;
            "LEFT_17_13": value  <= 0.46324449777603149414;
            "LEFT_17_14": value  <= 0.51322317123413085938;
            "LEFT_17_15": value  <= 0.66936898231506347656;
            "LEFT_17_16": value  <= 0.40538620948791498355;
            "LEFT_17_17": value  <= 0.64549958705902099609;
            "LEFT_17_18": value  <= 0.52704071998596191406;
            "LEFT_17_19": value  <= 0.38035470247268682309;
            "LEFT_17_20": value  <= 0.53394031524658203125;
            "LEFT_17_21": value  <= 0.35646161437034612485;
            "LEFT_17_22": value  <= 0.46719071269035339355;
            "LEFT_17_23": value  <= 0.51514732837677001953;
            "LEFT_17_24": value  <= 0.30416610836982732602;
            "LEFT_17_25": value  <= 0.64302957057952880859;
            "LEFT_17_26": value  <= 0.53074932098388671875;
            "LEFT_17_27": value  <= 0.46500471234321588687;
            "LEFT_17_28": value  <= 0.28496798872947687320;
            "LEFT_17_29": value  <= 0.29716458916664117984;
            "LEFT_17_30": value  <= 0.56310981512069702148;
            "LEFT_17_31": value  <= 0.44035780429840087891;
            "LEFT_17_32": value  <= 0.34210088849067687988;
            "LEFT_17_33": value  <= 0.46393430233001708984;
            "LEFT_17_34": value  <= 0.28201588988304138184;
            "LEFT_17_35": value  <= 0.52089059352874755859;
            "LEFT_17_36": value  <= 0.46637138724327087402;
            "LEFT_17_37": value  <= 0.52093499898910522461;
            "LEFT_17_38": value  <= 0.60631012916564941406;
            "LEFT_17_39": value  <= 0.46352049708366388492;
            "LEFT_17_40": value  <= 0.52894401550292968750;
            "LEFT_17_41": value  <= 0.77520018815994262695;
            "LEFT_17_42": value  <= 0.24280390143394470215;
            "LEFT_17_43": value  <= 0.57343649864196777344;
            "LEFT_17_44": value  <= 0.50298362970352172852;
            "LEFT_17_45": value  <= 0.60730451345443725586;
            "LEFT_17_46": value  <= 0.50152891874313354492;
            "LEFT_17_47": value  <= 0.66144287586212158203;
            "LEFT_17_48": value  <= 0.51808780431747436523;
            "LEFT_17_49": value  <= 0.47204169631004327945;
            "LEFT_17_50": value  <= 0.38050109148025512695;
            "LEFT_17_51": value  <= 0.29441660642623901367;
            "LEFT_17_52": value  <= 0.73461771011352539062;
            "LEFT_17_53": value  <= 0.54528760910034179688;
            "LEFT_17_54": value  <= 0.43988621234893798828;
            "LEFT_17_55": value  <= 0.47416868805885320493;
            "LEFT_17_56": value  <= 0.60445529222488403320;
            "LEFT_17_57": value  <= 0.24524590373039251157;
            "LEFT_17_58": value  <= 0.37328380346298217773;
            "LEFT_17_59": value  <= 0.54988098144531250000;
            "LEFT_17_60": value  <= 0.21399089694023129549;
            "LEFT_17_61": value  <= 0.46502870321273798160;
            "LEFT_17_62": value  <= 0.43874868750572210141;
            "LEFT_17_63": value  <= 0.52449727058410644531;
            "LEFT_17_64": value  <= 0.60568130016326904297;
            "LEFT_17_65": value  <= 0.20409290492534640227;
            "LEFT_17_66": value  <= 0.52376049757003784180;
            "LEFT_17_67": value  <= 0.49605339765548711606;
            "LEFT_17_68": value  <= 0.53513038158416748047;
            "LEFT_17_69": value  <= 0.46933668851852422543;
            "LEFT_17_70": value  <= 0.67913967370986938477;
            "LEFT_17_71": value  <= 0.36087390780448908023;
            "LEFT_17_72": value  <= 0.53000730276107788086;
            "LEFT_17_73": value  <= 0.51573169231414794922;
            "LEFT_17_74": value  <= 0.44104969501495361328;
            "LEFT_17_75": value  <= 0.54018551111221313477;
            "LEFT_17_76": value  <= 0.43682709336280822754;
            "LEFT_17_77": value  <= 0.42447990179061889648;
            "LEFT_17_78": value  <= 0.44969621300697332211;
            "LEFT_17_79": value  <= 0.52934932708740234375;
            "LEFT_17_80": value  <= 0.44832968711853027344;
            "LEFT_17_81": value  <= 0.45595070719718927554;
            "LEFT_17_82": value  <= 0.53417861461639404297;
            "LEFT_17_83": value  <= 0.56671887636184692383;
            "LEFT_17_84": value  <= 0.44212448596954351254;
            "LEFT_17_85": value  <= 0.42883709073066711426;
            "LEFT_17_86": value  <= 0.68995130062103271484;
            "LEFT_17_87": value  <= 0.22177790105342870541;
            "LEFT_17_88": value  <= 0.51362240314483642578;
            "LEFT_17_89": value  <= 0.48261928558349609375;
            "LEFT_17_90": value  <= 0.39228358864784240723;
            "LEFT_17_91": value  <= 0.50782018899917602539;
            "LEFT_17_92": value  <= 0.55204898118972778320;
            "LEFT_17_93": value  <= 0.39346051216125488281;
            "LEFT_17_94": value  <= 0.73706287145614624023;
            "LEFT_17_95": value  <= 0.51592797040939331055;
            "LEFT_17_96": value  <= 0.36728268861770629883;
            "LEFT_17_97": value  <= 0.50314939022064208984;
            "LEFT_17_98": value  <= 0.67675197124481201172;
            "LEFT_17_99": value  <= 0.52579981088638305664;
            "LEFT_17_100": value  <= 0.46962729096412658691;
            "LEFT_17_101": value  <= 0.43207129836082458496;
            "LEFT_17_102": value  <= 0.49977061152458190918;
            "LEFT_17_103": value  <= 0.42824178934097290039;
            "LEFT_17_104": value  <= 0.67721211910247802734;
            "LEFT_17_105": value  <= 0.53133970499038696289;
            "LEFT_17_106": value  <= 0.56600618362426757812;
            "LEFT_17_107": value  <= 0.37319138646125787906;
            "LEFT_17_108": value  <= 0.51899862289428710938;
            "LEFT_17_109": value  <= 0.29563739895820617676;
            "LEFT_17_110": value  <= 0.43471351265907287598;
            "LEFT_17_111": value  <= 0.32303300499916082211;
            "LEFT_17_112": value  <= 0.59754890203475952148;
            "LEFT_17_113": value  <= 0.47456780076026922055;
            "LEFT_17_114": value  <= 0.43244731426239008121;
            "LEFT_17_115": value  <= 0.15800529718399050627;
            "LEFT_17_116": value  <= 0.45176368951797490903;
            "LEFT_17_117": value  <= 0.41496479511260991879;
            "LEFT_17_118": value  <= 0.40390908718109130859;
            "LEFT_17_119": value  <= 0.47676518559455871582;
            "LEFT_17_120": value  <= 0.35862588882446289062;
            "LEFT_17_121": value  <= 0.47121399641036987305;
            "LEFT_17_122": value  <= 0.26610270142555242368;
            "LEFT_17_123": value  <= 0.51443397998809814453;
            "LEFT_17_124": value  <= 0.42849949002265930176;
            "LEFT_17_125": value  <= 0.38858351111412048340;
            "LEFT_17_126": value  <= 0.54125630855560302734;
            "LEFT_17_127": value  <= 0.48993051052093511410;
            "LEFT_17_128": value  <= 0.52867782115936279297;
            "LEFT_17_129": value  <= 0.60329902172088623047;
            "LEFT_17_130": value  <= 0.40844011306762700864;
            "LEFT_17_131": value  <= 0.48460629582405090332;
            "LEFT_17_132": value  <= 0.51647412776947021484;
            "LEFT_17_133": value  <= 0.56775820255279541016;
            "LEFT_17_134": value  <= 0.47314870357513427734;
            "LEFT_17_135": value  <= 0.52402430772781372070;
            "LEFT_17_136": value  <= 0.28370139002799987793;
            "LEFT_17_137": value  <= 0.74007177352905273438;
            "LEFT_17_138": value  <= 0.51191312074661254883;
            "LEFT_17_139": value  <= 0.49237880110740661621;
            "LEFT_17_140": value  <= 0.24347110092639920320;
            "LEFT_17_141": value  <= 0.59003108739852905273;
            "LEFT_17_142": value  <= 0.36473178863525390625;
            "LEFT_17_143": value  <= 0.60349482297897338867;
            "LEFT_17_144": value  <= 0.58189898729324340820;
            "LEFT_17_145": value  <= 0.52174758911132812500;
            "LEFT_17_146": value  <= 0.23607000708580019865;
            "LEFT_17_147": value  <= 0.64991867542266845703;
            "LEFT_17_148": value  <= 0.44133231043815607242;
            "LEFT_17_149": value  <= 0.43597310781478881836;
            "LEFT_17_150": value  <= 0.55040627717971801758;
            "LEFT_17_151": value  <= 0.40641129016876220703;
            "LEFT_17_152": value  <= 0.04735197126865389738;
            "LEFT_17_153": value  <= 0.48817330598831182309;
            "LEFT_17_154": value  <= 0.54000371694564819336;
            "LEFT_17_155": value  <= 0.48020479083061218262;
            "LEFT_17_156": value  <= 0.73877930641174316406;
            "LEFT_17_157": value  <= 0.52885460853576660156;
            "LEFT_17_158": value  <= 0.47508129477500921078;
            "LEFT_17_159": value  <= 0.38117301464080810547;
            "LEFT_18_0": value  <= 0.40191569924354547672;
            "LEFT_18_1": value  <= 0.33511489629745477847;
            "LEFT_18_2": value  <= 0.55577081441879272461;
            "LEFT_18_3": value  <= 0.42608588933944702148;
            "LEFT_18_4": value  <= 0.34942400455474847965;
            "LEFT_18_5": value  <= 0.40284991264343261719;
            "LEFT_18_6": value  <= 0.38069018721580510922;
            "LEFT_18_7": value  <= 0.26201000809669500180;
            "LEFT_18_8": value  <= 0.37997689843177800961;
            "LEFT_18_9": value  <= 0.44336450099945068359;
            "LEFT_18_10": value  <= 0.37196549773216247559;
            "LEFT_18_11": value  <= 0.55253958702087402344;
            "LEFT_18_12": value  <= 0.42645010352134710141;
            "LEFT_18_13": value  <= 0.43595260381698608398;
            "LEFT_18_14": value  <= 0.33901369571685791016;
            "LEFT_18_15": value  <= 0.45574560761451721191;
            "LEFT_18_16": value  <= 0.51348412036895751953;
            "LEFT_18_17": value  <= 0.39065781235694890805;
            "LEFT_18_18": value  <= 0.36796098947525018863;
            "LEFT_18_19": value  <= 0.72931021451950073242;
            "LEFT_18_20": value  <= 0.43453249335289001465;
            "LEFT_18_21": value  <= 0.25912800431251531430;
            "LEFT_18_22": value  <= 0.69222790002822875977;
            "LEFT_18_23": value  <= 0.53522628545761108398;
            "LEFT_18_24": value  <= 0.20405440032482149992;
            "LEFT_18_25": value  <= 0.68048888444900512695;
            "LEFT_18_26": value  <= 0.53106957674026489258;
            "LEFT_18_27": value  <= 0.57415628433227539062;
            "LEFT_18_28": value  <= 0.28317859768867492676;
            "LEFT_18_29": value  <= 0.33725079894065862485;
            "LEFT_18_30": value  <= 0.53066742420196533203;
            "LEFT_18_31": value  <= 0.54624962806701660156;
            "LEFT_18_32": value  <= 0.21578240394592290707;
            "LEFT_18_33": value  <= 0.64653122425079345703;
            "LEFT_18_34": value  <= 0.46176680922508239746;
            "LEFT_18_35": value  <= 0.52206891775131225586;
            "LEFT_18_36": value  <= 0.40145379304885858707;
            "LEFT_18_37": value  <= 0.47940391302108770200;
            "LEFT_18_38": value  <= 0.20341950654983520508;
            "LEFT_18_39": value  <= 0.76724731922149658203;
            "LEFT_18_40": value  <= 0.74903422594070434570;
            "LEFT_18_41": value  <= 0.53653037548065185547;
            "LEFT_18_42": value  <= 0.07401549816131590409;
            "LEFT_18_43": value  <= 0.28591030836105352231;
            "LEFT_18_44": value  <= 0.41916158795356750488;
            "LEFT_18_45": value  <= 0.62731927633285522461;
            "LEFT_18_46": value  <= 0.51599407196044921875;
            "LEFT_18_47": value  <= 0.58843767642974853516;
            "LEFT_18_48": value  <= 0.35605099797248840332;
            "LEFT_18_49": value  <= 0.59942889213562011719;
            "LEFT_18_50": value  <= 0.33454620838165277652;
            "LEFT_18_51": value  <= 0.55826562643051147461;
            "LEFT_18_52": value  <= 0.46236801147460937500;
            "LEFT_18_53": value  <= 0.65570747852325439453;
            "LEFT_18_54": value  <= 0.52695018053054809570;
            "LEFT_18_55": value  <= 0.46333730220794677734;
            "LEFT_18_56": value  <= 0.26896080374717712402;
            "LEFT_18_57": value  <= 0.54566031694412231445;
            "LEFT_18_58": value  <= 0.46489939093589782715;
            "LEFT_18_59": value  <= 0.53097039461135864258;
            "LEFT_18_60": value  <= 0.40747389197349548340;
            "LEFT_18_61": value  <= 0.19921760261058810149;
            "LEFT_18_62": value  <= 0.54385018348693847656;
            "LEFT_18_63": value  <= 0.42591789364814758301;
            "LEFT_18_64": value  <= 0.69041568040847778320;
            "LEFT_18_65": value  <= 0.45249149203300481625;
            "LEFT_18_66": value  <= 0.53703737258911132812;
            "LEFT_18_67": value  <= 0.64235579967498779297;
            "LEFT_18_68": value  <= 0.49884751439094537906;
            "LEFT_18_69": value  <= 0.54160261154174804688;
            "LEFT_18_70": value  <= 0.45763289928436279297;
            "LEFT_18_71": value  <= 0.53089731931686401367;
            "LEFT_18_72": value  <= 0.47056341171264648438;
            "LEFT_18_73": value  <= 0.44061261415481567383;
            "LEFT_18_74": value  <= 0.51290237903594970703;
            "LEFT_18_75": value  <= 0.31354710459709167480;
            "LEFT_18_76": value  <= 0.41193708777427667789;
            "LEFT_18_77": value  <= 0.61778062582015991211;
            "LEFT_18_78": value  <= 0.36543309688568120785;
            "LEFT_18_79": value  <= 0.34909150004386901855;
            "LEFT_18_80": value  <= 0.51662999391555786133;
            "LEFT_18_81": value  <= 0.50147360563278198242;
            "LEFT_18_82": value  <= 0.64707887172698974609;
            "LEFT_18_83": value  <= 0.32463788986206060239;
            "LEFT_18_84": value  <= 0.51919418573379516602;
            "LEFT_18_85": value  <= 0.49181339144706731625;
            "LEFT_18_86": value  <= 0.18368029594421389494;
            "LEFT_18_87": value  <= 0.52270537614822387695;
            "LEFT_18_88": value  <= 0.44902500510215759277;
            "LEFT_18_89": value  <= 0.48047870397567749023;
            "LEFT_18_90": value  <= 0.25210499763488769531;
            "LEFT_18_91": value  <= 0.59966957569122314453;
            "LEFT_18_92": value  <= 0.51537168025970458984;
            "LEFT_18_93": value  <= 0.66217190027236938477;
            "LEFT_18_94": value  <= 0.46333950757980352231;
            "LEFT_18_95": value  <= 0.36155730485916137695;
            "LEFT_18_96": value  <= 0.44428890943527221680;
            "LEFT_18_97": value  <= 0.51629352569580078125;
            "LEFT_18_98": value  <= 0.27896320819854741879;
            "LEFT_18_99": value  <= 0.49689841270446777344;
            "LEFT_18_100": value  <= 0.44456079602241521664;
            "LEFT_18_101": value  <= 0.02938820980489249834;
            "LEFT_18_102": value  <= 0.56993997097015380859;
            "LEFT_18_103": value  <= 0.43054661154747009277;
            "LEFT_18_104": value  <= 0.36803171038627630063;
            "LEFT_18_105": value  <= 0.48389169573783880063;
            "LEFT_18_106": value  <= 0.53252232074737548828;
            "LEFT_18_107": value  <= 0.48109480738639831543;
            "LEFT_18_108": value  <= 0.52002298831939697266;
            "LEFT_18_109": value  <= 0.49617099761962890625;
            "LEFT_18_110": value  <= 0.40602791309356689453;
            "LEFT_18_111": value  <= 0.46741139888763427734;
            "LEFT_18_112": value  <= 0.45191168785095220395;
            "LEFT_18_113": value  <= 0.28078991174697881528;
            "LEFT_18_114": value  <= 0.52955842018127441406;
            "LEFT_18_115": value  <= 0.54614001512527465820;
            "LEFT_18_116": value  <= 0.53291612863540649414;
            "LEFT_18_117": value  <= 0.45120179653167730160;
            "LEFT_18_118": value  <= 0.45778059959411621094;
            "LEFT_18_119": value  <= 0.52996039390563964844;
            "LEFT_18_120": value  <= 0.49590590596199041196;
            "LEFT_18_121": value  <= 0.51170790195465087891;
            "LEFT_18_122": value  <= 0.47363498806953430176;
            "LEFT_18_123": value  <= 0.52164179086685180664;
            "LEFT_18_124": value  <= 0.58098608255386352539;
            "LEFT_18_125": value  <= 0.53983622789382934570;
            "LEFT_18_126": value  <= 0.42492860555648798160;
            "LEFT_18_127": value  <= 0.52699637413024902344;
            "LEFT_18_128": value  <= 0.56330758333206176758;
            "LEFT_18_129": value  <= 0.53128892183303833008;
            "LEFT_18_130": value  <= 0.47017949819564819336;
            "LEFT_18_131": value  <= 0.00000000000000000000;
            "LEFT_18_132": value  <= 0.02374527975916860059;
            "LEFT_18_133": value  <= 0.31273230910301208496;
            "LEFT_18_134": value  <= 0.50090491771697998047;
            "LEFT_18_135": value  <= 0.63871437311172485352;
            "LEFT_18_136": value  <= 0.51368498802185058594;
            "LEFT_18_137": value  <= 0.55098438262939453125;
            "LEFT_18_138": value  <= 0.61623352766036987305;
            "LEFT_18_139": value  <= 0.61854577064514160156;
            "LEFT_18_140": value  <= 0.13826179504394531250;
            "LEFT_18_141": value  <= 0.46880578994750982114;
            "LEFT_18_142": value  <= 0.23685149848461151123;
            "LEFT_18_143": value  <= 0.58563941717147827148;
            "LEFT_18_144": value  <= 0.08690006285905839400;
            "LEFT_18_145": value  <= 0.51388370990753173828;
            "LEFT_18_146": value  <= 0.73536360263824462891;
            "LEFT_18_147": value  <= 0.38844060897827148438;
            "LEFT_18_148": value  <= 0.52234929800033569336;
            "LEFT_18_149": value  <= 0.49591061472892761230;
            "LEFT_18_150": value  <= 0.44448840618133550473;
            "LEFT_18_151": value  <= 0.53983712196350097656;
            "LEFT_18_152": value  <= 0.58542650938034057617;
            "LEFT_18_153": value  <= 0.46080690622329711914;
            "LEFT_18_154": value  <= 0.37911269068717962094;
            "LEFT_18_155": value  <= 0.59986090660095214844;
            "LEFT_18_156": value  <= 0.44842061400413507632;
            "LEFT_18_157": value  <= 0.54507470130920410156;
            "LEFT_18_158": value  <= 0.41182750463485717773;
            "LEFT_18_159": value  <= 0.57879078388214111328;
            "LEFT_18_160": value  <= 0.83978658914566040039;
            "LEFT_18_161": value  <= 0.24086110293865201082;
            "LEFT_18_162": value  <= 0.43553608655929570981;
            "LEFT_18_163": value  <= 0.54539710283279418945;
            "LEFT_18_164": value  <= 0.57710242271423339844;
            "LEFT_18_165": value  <= 0.51698678731918334961;
            "LEFT_18_166": value  <= 0.22032439708709719572;
            "LEFT_18_167": value  <= 0.50434082746505737305;
            "LEFT_18_168": value  <= 0.21862849593162539397;
            "LEFT_18_169": value  <= 0.50076818466186523438;
            "LEFT_18_170": value  <= 0.41298410296440130063;
            "LEFT_18_171": value  <= 0.54128682613372802734;
            "LEFT_18_172": value  <= 0.46055299043655401059;
            "LEFT_18_173": value  <= 0.52788549661636352539;
            "LEFT_18_174": value  <= 0.51296097040176391602;
            "LEFT_18_175": value  <= 0.48226919770240778140;
            "LEFT_18_176": value  <= 0.52483952045440673828;
            "LEFT_19_0": value  <= 0.34989839792251592465;
            "LEFT_19_1": value  <= 0.68166369199752807617;
            "LEFT_19_2": value  <= 0.55857062339782714844;
            "LEFT_19_3": value  <= 0.53650361299514770508;
            "LEFT_19_4": value  <= 0.36390951275825500488;
            "LEFT_19_5": value  <= 0.28591570258140558414;
            "LEFT_19_6": value  <= 0.52365237474441528320;
            "LEFT_19_7": value  <= 0.47503221035003662109;
            "LEFT_19_8": value  <= 0.33433759212493902035;
            "LEFT_19_9": value  <= 0.51921808719635009766;
            "LEFT_19_10": value  <= 0.29298439621925348453;
            "LEFT_19_11": value  <= 0.36868458986282348633;
            "LEFT_19_12": value  <= 0.36321839690208440610;
            "LEFT_19_13": value  <= 0.58706837892532348633;
            "LEFT_19_14": value  <= 0.31958949565887451172;
            "LEFT_19_15": value  <= 0.63018590211868286133;
            "LEFT_19_16": value  <= 0.19770480692386629973;
            "LEFT_19_17": value  <= 0.49541321396827697754;
            "LEFT_19_18": value  <= 0.51644277572631835938;
            "LEFT_19_19": value  <= 0.23152460157871249113;
            "LEFT_19_20": value  <= 0.46642971038818359375;
            "LEFT_19_21": value  <= 0.52208751440048217773;
            "LEFT_19_22": value  <= 0.50792771577835083008;
            "LEFT_19_23": value  <= 0.48859509825706481934;
            "LEFT_19_24": value  <= 0.51972568035125732422;
            "LEFT_19_25": value  <= 0.61534678936004638672;
            "LEFT_19_26": value  <= 0.26373448967933660336;
            "LEFT_19_27": value  <= 0.22875219583511349764;
            "LEFT_19_28": value  <= 0.69533038139343261719;
            "LEFT_19_29": value  <= 0.54506552219390869141;
            "LEFT_19_30": value  <= 0.60913878679275512695;
            "LEFT_19_31": value  <= 0.52410632371902465820;
            "LEFT_19_32": value  <= 0.53879290819168090820;
            "LEFT_19_33": value  <= 0.42926910519599920102;
            "LEFT_19_34": value  <= 0.37923479080200200864;
            "LEFT_19_35": value  <= 0.52372831106185913086;
            "LEFT_19_36": value  <= 0.19476559758186340332;
            "LEFT_19_37": value  <= 0.60112851858139038086;
            "LEFT_19_38": value  <= 0.50097537040710449219;
            "LEFT_19_39": value  <= 0.48621898889541631528;
            "LEFT_19_40": value  <= 0.50002187490463256836;
            "LEFT_19_41": value  <= 0.55301171541213989258;
            "LEFT_19_42": value  <= 0.41786059737205510922;
            "LEFT_19_43": value  <= 0.49971699714660650082;
            "LEFT_19_44": value  <= 0.53318071365356445312;
            "LEFT_19_45": value  <= 0.57559251785278320312;
            "LEFT_19_46": value  <= 0.45769768953323358707;
            "LEFT_19_47": value  <= 0.43803969025611877441;
            "LEFT_19_48": value  <= 0.51630318164825439453;
            "LEFT_19_49": value  <= 0.60729467868804931641;
            "LEFT_19_50": value  <= 0.32924759387969970703;
            "LEFT_19_51": value  <= 0.48297679424285888672;
            "LEFT_19_52": value  <= 0.46606799960136408023;
            "LEFT_19_53": value  <= 0.52048492431640625000;
            "LEFT_19_54": value  <= 0.51673221588134765625;
            "LEFT_19_55": value  <= 0.64064931869506835938;
            "LEFT_19_56": value  <= 0.58972930908203125000;
            "LEFT_19_57": value  <= 0.54415607452392578125;
            "LEFT_19_58": value  <= 0.21431629359722140227;
            "LEFT_19_59": value  <= 0.53864240646362304688;
            "LEFT_19_60": value  <= 0.57511842250823974609;
            "LEFT_19_61": value  <= 0.54219377040863037109;
            "LEFT_19_62": value  <= 0.40779209136962890625;
            "LEFT_19_63": value  <= 0.42292758822441101074;
            "LEFT_19_64": value  <= 0.65963757038116455078;
            "LEFT_19_65": value  <= 0.42511358857154851743;
            "LEFT_19_66": value  <= 0.52592468261718750000;
            "LEFT_19_67": value  <= 0.46717229485511779785;
            "LEFT_19_68": value  <= 0.57110661268234252930;
            "LEFT_19_69": value  <= 0.52641981840133666992;
            "LEFT_19_70": value  <= 0.38917380571365361996;
            "LEFT_19_71": value  <= 0.57958728075027465820;
            "LEFT_19_72": value  <= 0.23776030540466311369;
            "LEFT_19_73": value  <= 0.48766261339187622070;
            "LEFT_19_74": value  <= 0.51680880784988403320;
            "LEFT_19_75": value  <= 0.54466491937637329102;
            "LEFT_19_76": value  <= 0.46878978610038757324;
            "LEFT_19_77": value  <= 0.51934438943862915039;
            "LEFT_19_78": value  <= 0.49717310070991521664;
            "LEFT_19_79": value  <= 0.51659947633743286133;
            "LEFT_19_80": value  <= 0.40584719181060791016;
            "LEFT_19_81": value  <= 0.34450569748878479004;
            "LEFT_19_82": value  <= 0.45948630571365361996;
            "LEFT_19_83": value  <= 0.16804009675979608707;
            "LEFT_19_84": value  <= 0.38615968823432922363;
            "LEFT_19_85": value  <= 0.55179792642593383789;
            "LEFT_19_86": value  <= 0.79994601011276245117;
            "LEFT_19_87": value  <= 0.40859758853912347965;
            "LEFT_19_88": value  <= 0.54704052209854125977;
            "LEFT_19_89": value  <= 0.49889969825744628906;
            "LEFT_19_90": value  <= 0.67536902427673339844;
            "LEFT_19_91": value  <= 0.54158538579940795898;
            "LEFT_19_92": value  <= 0.22585099935531618986;
            "LEFT_19_93": value  <= 0.62565547227859497070;
            "LEFT_19_94": value  <= 0.39477849006652832031;
            "LEFT_19_95": value  <= 0.47525110840797418765;
            "LEFT_19_96": value  <= 0.60411047935485839844;
            "LEFT_19_97": value  <= 0.42582759261131292172;
            "LEFT_19_98": value  <= 0.52334201335906982422;
            "LEFT_19_99": value  <= 0.63718891143798828125;
            "LEFT_19_100": value  <= 0.53747057914733886719;
            "LEFT_19_101": value  <= 0.46387958526611328125;
            "LEFT_19_102": value  <= 0.46886560320854192563;
            "LEFT_19_103": value  <= 0.52043187618255615234;
            "LEFT_19_104": value  <= 0.16303719580173489656;
            "LEFT_19_105": value  <= 0.57744592428207397461;
            "LEFT_19_106": value  <= 0.39771759510040277652;
            "LEFT_19_107": value  <= 0.60465282201766967773;
            "LEFT_19_108": value  <= 0.39967238903045648746;
            "LEFT_19_109": value  <= 0.47121581435203552246;
            "LEFT_19_110": value  <= 0.41095849871635442563;
            "LEFT_19_111": value  <= 0.52029937505722045898;
            "LEFT_19_112": value  <= 0.65666097402572631836;
            "LEFT_19_113": value  <= 0.51286739110946655273;
            "LEFT_19_114": value  <= 0.65807867050170898438;
            "LEFT_19_115": value  <= 0.51464450359344482422;
            "LEFT_19_116": value  <= 0.38366019725799560547;
            "LEFT_19_117": value  <= 0.50855928659439086914;
            "LEFT_19_118": value  <= 0.51387631893157958984;
            "LEFT_19_119": value  <= 0.59896552562713623047;
            "LEFT_19_120": value  <= 0.45094868540763860532;
            "LEFT_19_121": value  <= 0.34967708587646478824;
            "LEFT_19_122": value  <= 0.11205369979143139925;
            "LEFT_19_123": value  <= 0.51481968164443969727;
            "LEFT_19_124": value  <= 0.40849998593330377750;
            "LEFT_19_125": value  <= 0.63941049575805664062;
            "LEFT_19_126": value  <= 0.47075539827346801758;
            "LEFT_19_127": value  <= 0.45413690805435180664;
            "LEFT_19_128": value  <= 0.43339619040489202328;
            "LEFT_19_129": value  <= 0.45796871185302728824;
            "LEFT_19_130": value  <= 0.43246439099311828613;
            "LEFT_19_131": value  <= 0.52572208642959594727;
            "LEFT_19_132": value  <= 0.60430181026458740234;
            "LEFT_19_133": value  <= 0.45982548594474792480;
            "LEFT_19_134": value  <= 0.41307520866394037418;
            "LEFT_19_135": value  <= 0.40430399775505071469;
            "LEFT_19_136": value  <= 0.44949638843536382504;
            "LEFT_19_137": value  <= 0.51775109767913818359;
            "LEFT_19_138": value  <= 0.19880190491676330566;
            "LEFT_19_139": value  <= 0.66447502374649047852;
            "LEFT_19_140": value  <= 0.38983049988746637515;
            "LEFT_19_141": value  <= 0.48018088936805730649;
            "LEFT_19_142": value  <= 0.52109199762344360352;
            "LEFT_19_143": value  <= 0.61545419692993164062;
            "LEFT_19_144": value  <= 0.39759421348571777344;
            "LEFT_19_145": value  <= 0.49791380763053888492;
            "LEFT_19_146": value  <= 0.49844971299171447754;
            "LEFT_19_147": value  <= 0.59049648046493530273;
            "LEFT_19_148": value  <= 0.41995579004287719727;
            "LEFT_19_149": value  <= 0.54186028242111206055;
            "LEFT_19_150": value  <= 0.37259390950202941895;
            "LEFT_19_151": value  <= 0.64789611101150512695;
            "LEFT_19_152": value  <= 0.46823391318321228027;
            "LEFT_19_153": value  <= 0.54585301876068115234;
            "LEFT_19_154": value  <= 0.36901599168777471371;
            "LEFT_19_155": value  <= 0.60505628585815429688;
            "LEFT_19_156": value  <= 0.20170800387859338931;
            "LEFT_19_157": value  <= 0.57131487131118774414;
            "LEFT_19_158": value  <= 0.42153888940811157227;
            "LEFT_19_159": value  <= 0.51361519098281860352;
            "LEFT_19_160": value  <= 0.70273578166961669922;
            "LEFT_19_161": value  <= 0.43174090981483459473;
            "LEFT_19_162": value  <= 0.59426987171173095703;
            "LEFT_19_163": value  <= 0.61915689706802368164;
            "LEFT_19_164": value  <= 0.52566647529602050781;
            "LEFT_19_165": value  <= 0.52378678321838378906;
            "LEFT_19_166": value  <= 0.21304459869861600008;
            "LEFT_19_167": value  <= 0.48140418529510498047;
            "LEFT_19_168": value  <= 0.64825797080993652344;
            "LEFT_19_169": value  <= 0.45819279551506042480;
            "LEFT_19_170": value  <= 0.52320867776870727539;
            "LEFT_19_171": value  <= 0.55562019348144531250;
            "LEFT_19_172": value  <= 0.52294427156448364258;
            "LEFT_19_173": value  <= 0.62986820936203002930;
            "LEFT_19_174": value  <= 0.72282809019088745117;
            "LEFT_19_175": value  <= 0.22695130109786990080;
            "LEFT_19_176": value  <= 0.52370971441268920898;
            "LEFT_19_177": value  <= 0.47737509012222290039;
            "LEFT_19_178": value  <= 0.71469759941101074219;
            "LEFT_19_179": value  <= 0.26352968811988830566;
            "LEFT_19_180": value  <= 0.36237570643424987793;
            "LEFT_19_181": value  <= 0.47059321403503417969;
            "LEFT_20_0": value  <= 0.38605189323425287418;
            "LEFT_20_1": value  <= 0.43856549263000488281;
            "LEFT_20_2": value  <= 0.54871010780334472656;
            "LEFT_20_3": value  <= 0.32305321097373962402;
            "LEFT_20_4": value  <= 0.50916397571563720703;
            "LEFT_20_5": value  <= 0.41781538724899291992;
            "LEFT_20_6": value  <= 0.28991821408271789551;
            "LEFT_20_7": value  <= 0.42801249027252197266;
            "LEFT_20_8": value  <= 0.40448719263076782227;
            "LEFT_20_9": value  <= 0.42717689275741582700;
            "LEFT_20_10": value  <= 0.39627239108085632324;
            "LEFT_20_11": value  <= 0.47271779179573059082;
            "LEFT_20_12": value  <= 0.56030082702636718750;
            "LEFT_20_13": value  <= 0.52259171009063720703;
            "LEFT_20_14": value  <= 0.39990758895874017886;
            "LEFT_20_15": value  <= 0.46783858537673950195;
            "LEFT_20_16": value  <= 0.34939670562744140625;
            "LEFT_20_17": value  <= 0.61858189105987548828;
            "LEFT_20_18": value  <= 0.52853411436080932617;
            "LEFT_20_19": value  <= 0.53606408834457397461;
            "LEFT_20_20": value  <= 0.45582920312881469727;
            "LEFT_20_21": value  <= 0.36802300810813898257;
            "LEFT_20_22": value  <= 0.39605951309204101562;
            "LEFT_20_23": value  <= 0.70204448699951171875;
            "LEFT_20_24": value  <= 0.50491642951965332031;
            "LEFT_20_25": value  <= 0.26726329326629638672;
            "LEFT_20_26": value  <= 0.45794829726219177246;
            "LEFT_20_27": value  <= 0.31715941429138178043;
            "LEFT_20_28": value  <= 0.52653628587722778320;
            "LEFT_20_29": value  <= 0.53324568271636962891;
            "LEFT_20_30": value  <= 0.45933109521865850278;
            "LEFT_20_31": value  <= 0.44379639625549321957;
            "LEFT_20_32": value  <= 0.46803238987922668457;
            "LEFT_20_33": value  <= 0.37096318602561950684;
            "LEFT_20_34": value  <= 0.47235551476478582211;
            "LEFT_20_35": value  <= 0.44923940300941467285;
            "LEFT_20_36": value  <= 0.44068640470504760742;
            "LEFT_20_37": value  <= 0.46824169158935552426;
            "LEFT_20_38": value  <= 0.50793921947479248047;
            "LEFT_20_39": value  <= 0.56010371446609497070;
            "LEFT_20_40": value  <= 0.22075350582599639893;
            "LEFT_20_41": value  <= 0.65312159061431884766;
            "LEFT_20_42": value  <= 0.49679630994796747379;
            "LEFT_20_43": value  <= 0.48989468812942510434;
            "LEFT_20_44": value  <= 0.39271169900894170590;
            "LEFT_20_45": value  <= 0.56133252382278442383;
            "LEFT_20_46": value  <= 0.44728800654411321469;
            "LEFT_20_47": value  <= 0.38405328989028930664;
            "LEFT_20_48": value  <= 0.58439838886260986328;
            "LEFT_20_49": value  <= 0.54392218589782714844;
            "LEFT_20_50": value  <= 0.12884649634361269865;
            "LEFT_20_51": value  <= 0.49512979388236999512;
            "LEFT_20_52": value  <= 0.39465999603271478824;
            "LEFT_20_53": value  <= 0.48975038528442377261;
            "LEFT_20_54": value  <= 0.32454401254653930664;
            "LEFT_20_55": value  <= 0.15819530189037320222;
            "LEFT_20_56": value  <= 0.46809351444244390317;
            "LEFT_20_57": value  <= 0.52116978168487548828;
            "LEFT_20_58": value  <= 0.57683861255645751953;
            "LEFT_20_59": value  <= 0.45077630877494812012;
            "LEFT_20_60": value  <= 0.54608201980590820312;
            "LEFT_20_61": value  <= 0.53718560934066772461;
            "LEFT_20_62": value  <= 0.44712871313095092773;
            "LEFT_20_63": value  <= 0.44993931055068969727;
            "LEFT_20_64": value  <= 0.55161732435226440430;
            "LEFT_20_65": value  <= 0.51941901445388793945;
            "LEFT_20_66": value  <= 0.38307058811187738590;
            "LEFT_20_67": value  <= 0.48910909891128540039;
            "LEFT_20_68": value  <= 0.74136817455291748047;
            "LEFT_20_69": value  <= 0.36488190293312072754;
            "LEFT_20_70": value  <= 0.51004928350448608398;
            "LEFT_20_71": value  <= 0.52324420213699340820;
            "LEFT_20_72": value  <= 0.46481490135192871094;
            "LEFT_20_73": value  <= 0.59303098917007446289;
            "LEFT_20_74": value  <= 0.38704779744148248843;
            "LEFT_20_75": value  <= 0.55225032567977905273;
            "LEFT_20_76": value  <= 0.45462208986282348633;
            "LEFT_20_77": value  <= 0.53457391262054443359;
            "LEFT_20_78": value  <= 0.39678159356117248535;
            "LEFT_20_79": value  <= 0.28296428918838500977;
            "LEFT_20_80": value  <= 0.45900669693946838379;
            "LEFT_20_81": value  <= 0.52314108610153198242;
            "LEFT_20_82": value  <= 0.43972569704055791684;
            "LEFT_20_83": value  <= 0.31350791454315191098;
            "LEFT_20_84": value  <= 0.32132729887962341309;
            "LEFT_20_85": value  <= 0.63875448703765869141;
            "LEFT_20_86": value  <= 0.27591320872306818179;
            "LEFT_20_87": value  <= 0.46856409311294561215;
            "LEFT_20_88": value  <= 0.51752072572708129883;
            "LEFT_20_89": value  <= 0.20691369473934170808;
            "LEFT_20_90": value  <= 0.61340910196304321289;
            "LEFT_20_91": value  <= 0.54541081190109252930;
            "LEFT_20_92": value  <= 0.63444852828979492188;
            "LEFT_20_93": value  <= 0.52926832437515258789;
            "LEFT_20_94": value  <= 0.43929880857467651367;
            "LEFT_20_95": value  <= 0.58988320827484130859;
            "LEFT_20_96": value  <= 0.40693649649620061703;
            "LEFT_20_97": value  <= 0.51827257871627807617;
            "LEFT_20_98": value  <= 0.13075779378414151277;
            "LEFT_20_99": value  <= 0.64210057258605957031;
            "LEFT_20_100": value  <= 0.04776934906840320239;
            "LEFT_20_101": value  <= 0.46162670850753778629;
            "LEFT_20_102": value  <= 0.62618541717529296875;
            "LEFT_20_103": value  <= 0.53844177722930908203;
            "LEFT_20_104": value  <= 0.38040471076965332031;
            "LEFT_20_105": value  <= 0.45543101429939270020;
            "LEFT_20_106": value  <= 0.65969580411911010742;
            "LEFT_20_107": value  <= 0.51954662799835205078;
            "LEFT_20_108": value  <= 0.52291762828826904297;
            "LEFT_20_109": value  <= 0.63528877496719360352;
            "LEFT_20_110": value  <= 0.38245460391044622250;
            "LEFT_20_111": value  <= 0.49504399299621582031;
            "LEFT_20_112": value  <= 0.49523359537124628238;
            "LEFT_20_113": value  <= 0.75427287817001342773;
            "LEFT_20_114": value  <= 0.36993029713630681821;
            "LEFT_20_115": value  <= 0.66891789436340332031;
            "LEFT_20_116": value  <= 0.49833008646965032407;
            "LEFT_20_117": value  <= 0.45744240283966058902;
            "LEFT_20_118": value  <= 0.51317447423934936523;
            "LEFT_20_119": value  <= 0.43617001175880432129;
            "LEFT_20_120": value  <= 0.46827208995819091797;
            "LEFT_20_121": value  <= 0.43292450904846191406;
            "LEFT_20_122": value  <= 0.53700572252273559570;
            "LEFT_20_123": value  <= 0.51372742652893066406;
            "LEFT_20_124": value  <= 0.41120609641075128726;
            "LEFT_20_125": value  <= 0.54046237468719482422;
            "LEFT_20_126": value  <= 0.43559691309928888492;
            "LEFT_20_127": value  <= 0.59951752424240112305;
            "LEFT_20_128": value  <= 0.49502879381179809570;
            "LEFT_20_129": value  <= 0.63972991704940795898;
            "LEFT_20_130": value  <= 0.10016699880361559782;
            "LEFT_20_131": value  <= 0.33123299479484558105;
            "LEFT_20_132": value  <= 0.44063639640808111020;
            "LEFT_20_133": value  <= 0.27995899319648742676;
            "LEFT_20_134": value  <= 0.69875800609588623047;
            "LEFT_20_135": value  <= 0.49832889437675481625;
            "LEFT_20_136": value  <= 0.29823330044746398926;
            "LEFT_20_137": value  <= 0.53084421157836914062;
            "LEFT_20_138": value  <= 0.20379640161991119385;
            "LEFT_20_139": value  <= 0.50256967544555664062;
            "LEFT_20_140": value  <= 0.49600529670715332031;
            "LEFT_20_141": value  <= 0.56030637025833129883;
            "LEFT_20_142": value  <= 0.52055621147155761719;
            "LEFT_20_143": value  <= 0.52216529846191406250;
            "LEFT_20_144": value  <= 0.60226827859878540039;
            "LEFT_20_145": value  <= 0.40704470872879028320;
            "LEFT_20_146": value  <= 0.46018350124359130859;
            "LEFT_20_147": value  <= 0.53982520103454589844;
            "LEFT_20_148": value  <= 0.52015632390975952148;
            "LEFT_20_149": value  <= 0.46423879265785217285;
            "LEFT_20_150": value  <= 0.61985671520233154297;
            "LEFT_20_151": value  <= 0.68373328447341918945;
            "LEFT_20_152": value  <= 0.43448030948638921567;
            "LEFT_20_153": value  <= 0.47600790858268737793;
            "LEFT_20_154": value  <= 0.50909858942031860352;
            "LEFT_20_155": value  <= 0.55700647830963134766;
            "LEFT_20_156": value  <= 0.53568458557128906250;
            "LEFT_20_157": value  <= 0.44398030638694757632;
            "LEFT_20_158": value  <= 0.40422949194908142090;
            "LEFT_20_159": value  <= 0.49276518821716308594;
            "LEFT_20_160": value  <= 0.80062937736511230469;
            "LEFT_20_161": value  <= 0.39460548758506780453;
            "LEFT_20_162": value  <= 0.02132499031722550134;
            "LEFT_20_163": value  <= 0.40127959847450261899;
            "LEFT_20_164": value  <= 0.46424189209938049316;
            "LEFT_20_165": value  <= 0.65021592378616333008;
            "LEFT_20_166": value  <= 0.52647089958190917969;
            "LEFT_20_167": value  <= 0.48791998624801641293;
            "LEFT_20_168": value  <= 0.39172801375389099121;
            "LEFT_20_169": value  <= 0.58375990390777587891;
            "LEFT_20_170": value  <= 0.12619839608669281006;
            "LEFT_20_171": value  <= 0.57225137948989868164;
            "LEFT_20_172": value  <= 0.52732622623443603516;
            "LEFT_20_173": value  <= 0.44500669836997991391;
            "LEFT_20_174": value  <= 0.57576531171798706055;
            "LEFT_20_175": value  <= 0.18843810260295870695;
            "LEFT_20_176": value  <= 0.65897899866104125977;
            "LEFT_20_177": value  <= 0.52594298124313354492;
            "LEFT_20_178": value  <= 0.53552711009979248047;
            "LEFT_20_179": value  <= 0.50344067811965942383;
            "LEFT_20_180": value  <= 0.47566050291061401367;
            "LEFT_20_181": value  <= 0.53696119785308837891;
            "LEFT_20_182": value  <= 0.49686419963836669922;
            "LEFT_20_183": value  <= 0.49307331442832952328;
            "LEFT_20_184": value  <= 0.52052050828933715820;
            "LEFT_20_185": value  <= 0.54835551977157592773;
            "LEFT_20_186": value  <= 0.46899020671844482422;
            "LEFT_20_187": value  <= 0.51711422204971313477;
            "LEFT_20_188": value  <= 0.52199780941009521484;
            "LEFT_20_189": value  <= 0.58603698015213012695;
            "LEFT_20_190": value  <= 0.17492769658565521240;
            "LEFT_20_191": value  <= 0.43425890803337102719;
            "LEFT_20_192": value  <= 0.47651869058609008789;
            "LEFT_20_193": value  <= 0.52621912956237792969;
            "LEFT_20_194": value  <= 0.48040691018104547672;
            "LEFT_20_195": value  <= 0.41208469867706298828;
            "LEFT_20_196": value  <= 0.47403728961944580078;
            "LEFT_20_197": value  <= 0.24687920510768890381;
            "LEFT_20_198": value  <= 0.57562941312789916992;
            "LEFT_20_199": value  <= 0.51696258783340454102;
            "LEFT_20_200": value  <= 0.38720148801803588867;
            "LEFT_20_201": value  <= 0.48530489206314092465;
            "LEFT_20_202": value  <= 0.51173150539398193359;
            "LEFT_20_203": value  <= 0.56927400827407836914;
            "LEFT_20_204": value  <= 0.25560128688812261410;
            "LEFT_20_205": value  <= 0.48108729720115661621;
            "LEFT_20_206": value  <= 0.49711948633193969727;
            "LEFT_20_207": value  <= 0.49400109052658081055;
            "LEFT_20_208": value  <= 0.50076121091842651367;
            "LEFT_20_209": value  <= 0.70595788955688476562;
            "LEFT_20_210": value  <= 0.51286202669143676758;
            "LEFT_21_0": value  <= 0.64707571268081665039;
            "LEFT_21_1": value  <= 0.39998221397399902344;
            "LEFT_21_2": value  <= 0.35587701201438898257;
            "LEFT_21_3": value  <= 0.42565348744392400571;
            "LEFT_21_4": value  <= 0.36829081177711492368;
            "LEFT_21_5": value  <= 0.54524701833724975586;
            "LEFT_21_6": value  <= 0.52390581369400024414;
            "LEFT_21_7": value  <= 0.43206891417503362485;
            "LEFT_21_8": value  <= 0.45046371221542358398;
            "LEFT_21_9": value  <= 0.43134251236915588379;
            "LEFT_21_10": value  <= 0.53266030550003051758;
            "LEFT_21_11": value  <= 0.43051639199256902524;
            "LEFT_21_12": value  <= 0.42359709739685058594;
            "LEFT_21_13": value  <= 0.53030598163604736328;
            "LEFT_21_14": value  <= 0.35571089386940002441;
            "LEFT_21_15": value  <= 0.52253627777099609375;
            "LEFT_21_16": value  <= 0.36241859197616582700;
            "LEFT_21_17": value  <= 0.54744768142700195312;
            "LEFT_21_18": value  <= 0.37404221296310430356;
            "LEFT_21_19": value  <= 0.58930522203445434570;
            "LEFT_21_20": value  <= 0.40845820307731628418;
            "LEFT_21_21": value  <= 0.37774550914764398746;
            "LEFT_21_22": value  <= 0.29636120796203607730;
            "LEFT_21_23": value  <= 0.48776328563690191098;
            "LEFT_21_24": value  <= 0.43669110536575317383;
            "LEFT_21_25": value  <= 0.31281578540802001953;
            "LEFT_21_26": value  <= 0.65602248907089233398;
            "LEFT_21_27": value  <= 0.51726800203323364258;
            "LEFT_21_28": value  <= 0.40844461321830749512;
            "LEFT_21_29": value  <= 0.49669221043586730957;
            "LEFT_21_30": value  <= 0.59082370996475219727;
            "LEFT_21_31": value  <= 0.53151607513427734375;
            "LEFT_21_32": value  <= 0.23340409994125368986;
            "LEFT_21_33": value  <= 0.58809357881546020508;
            "LEFT_21_34": value  <= 0.49837771058082580566;
            "LEFT_21_35": value  <= 0.58721381425857543945;
            "LEFT_21_36": value  <= 0.51311892271041870117;
            "LEFT_21_37": value  <= 0.53393721580505371094;
            "LEFT_21_38": value  <= 0.43133831024169921875;
            "LEFT_21_39": value  <= 0.26753368973732000180;
            "LEFT_21_40": value  <= 0.49738699197769170590;
            "LEFT_21_41": value  <= 0.55297082662582397461;
            "LEFT_21_42": value  <= 0.56295841932296752930;
            "LEFT_21_43": value  <= 0.67062127590179443359;
            "LEFT_21_44": value  <= 0.52394217252731323242;
            "LEFT_21_45": value  <= 0.47994381189346307925;
            "LEFT_21_46": value  <= 0.69300097227096557617;
            "LEFT_21_47": value  <= 0.40996238589286798648;
            "LEFT_21_48": value  <= 0.32834759354591369629;
            "LEFT_21_49": value  <= 0.49780470132827758789;
            "LEFT_21_50": value  <= 0.46611601114273071289;
            "LEFT_21_51": value  <= 0.23346449434757229890;
            "LEFT_21_52": value  <= 0.11836539953947070036;
            "LEFT_21_53": value  <= 0.53250199556350708008;
            "LEFT_21_54": value  <= 0.62787622213363647461;
            "LEFT_21_55": value  <= 0.34034150838851928711;
            "LEFT_21_56": value  <= 0.36104118824005132504;
            "LEFT_21_57": value  <= 0.48842659592628479004;
            "LEFT_21_58": value  <= 0.26259300112724298648;
            "LEFT_21_59": value  <= 0.43407949805259710141;
            "LEFT_21_60": value  <= 0.65079987049102783203;
            "LEFT_21_61": value  <= 0.38265028595924377441;
            "LEFT_21_62": value  <= 0.32333680987358087711;
            "LEFT_21_63": value  <= 0.51776039600372314453;
            "LEFT_21_64": value  <= 0.40208509564399719238;
            "LEFT_21_65": value  <= 0.63150721788406372070;
            "LEFT_21_66": value  <= 0.47024598717689508609;
            "LEFT_21_67": value  <= 0.36503839492797851562;
            "LEFT_21_68": value  <= 0.51661008596420288086;
            "LEFT_21_69": value  <= 0.73758941888809204102;
            "LEFT_21_70": value  <= 0.44232261180877691098;
            "LEFT_21_71": value  <= 0.59763962030410766602;
            "LEFT_21_72": value  <= 0.59559392929077148438;
            "LEFT_21_73": value  <= 0.53498882055282592773;
            "LEFT_21_74": value  <= 0.50491911172866821289;
            "LEFT_21_75": value  <= 0.25501778721809392758;
            "LEFT_21_76": value  <= 0.44248610734939580746;
            "LEFT_21_77": value  <= 0.53195142745971679688;
            "LEFT_21_78": value  <= 0.40876591205596918277;
            "LEFT_21_79": value  <= 0.56745791435241699219;
            "LEFT_21_80": value  <= 0.41294258832931518555;
            "LEFT_21_81": value  <= 0.50601941347122192383;
            "LEFT_21_82": value  <= 0.59796321392059326172;
            "LEFT_21_83": value  <= 0.41743651032447820493;
            "LEFT_21_84": value  <= 0.56158047914505004883;
            "LEFT_21_85": value  <= 0.40761870145797729492;
            "LEFT_21_86": value  <= 0.43472939729690551758;
            "LEFT_21_87": value  <= 0.16593049466609960385;
            "LEFT_21_88": value  <= 0.49618190526962280273;
            "LEFT_21_89": value  <= 0.48682639002799987793;
            "LEFT_21_90": value  <= 0.62843251228332519531;
            "LEFT_21_91": value  <= 0.55750000476837158203;
            "LEFT_21_92": value  <= 0.41157621145248407535;
            "LEFT_21_93": value  <= 0.47300729155540471860;
            "LEFT_21_94": value  <= 0.49718868732452392578;
            "LEFT_21_95": value  <= 0.53721177577972412109;
            "LEFT_21_96": value  <= 0.53668838739395141602;
            "LEFT_21_97": value  <= 0.34355181455612182617;
            "LEFT_21_98": value  <= 0.47667920589447021484;
            "LEFT_21_99": value  <= 0.50293159484863281250;
            "LEFT_21_100": value  <= 0.40160921216011047363;
            "LEFT_21_101": value  <= 0.40883159637451171875;
            "LEFT_21_102": value  <= 0.40756770968437200375;
            "LEFT_21_103": value  <= 0.49132829904556268863;
            "LEFT_21_104": value  <= 0.50316721200942993164;
            "LEFT_21_105": value  <= 0.49497890472412109375;
            "LEFT_21_106": value  <= 0.53283667564392089844;
            "LEFT_21_107": value  <= 0.49915251135826110840;
            "LEFT_21_108": value  <= 0.45735040307044977359;
            "LEFT_21_109": value  <= 0.46043589711189270020;
            "LEFT_21_110": value  <= 0.39693889021873468570;
            "LEFT_21_111": value  <= 0.58083200454711914062;
            "LEFT_21_112": value  <= 0.43512108922004699707;
            "LEFT_21_113": value  <= 0.53550601005554199219;
            "LEFT_21_114": value  <= 0.50181388854980468750;
            "LEFT_21_115": value  <= 0.12250760197639469495;
            "LEFT_21_116": value  <= 0.47317668795585632324;
            "LEFT_21_117": value  <= 0.54305320978164672852;
            "LEFT_21_118": value  <= 0.40310400724411010742;
            "LEFT_21_119": value  <= 0.43081268668174738101;
            "LEFT_21_120": value  <= 0.62198299169540405273;
            "LEFT_21_121": value  <= 0.53793638944625854492;
            "LEFT_21_122": value  <= 0.52816402912139892578;
            "LEFT_21_123": value  <= 0.25820928812026977539;
            "LEFT_21_124": value  <= 0.47786930203437810727;
            "LEFT_21_125": value  <= 0.53409922122955322266;
            "LEFT_21_126": value  <= 0.49657610058784490414;
            "LEFT_21_127": value  <= 0.64149940013885498047;
            "LEFT_21_128": value  <= 0.45223200321197509766;
            "LEFT_21_129": value  <= 0.27647489309310907535;
            "LEFT_21_130": value  <= 0.51419419050216674805;
            "LEFT_21_131": value  <= 0.50606489181518554688;
            "LEFT_21_132": value  <= 0.51953881978988647461;
            "LEFT_21_133": value  <= 0.49623650312423711606;
            "LEFT_21_134": value  <= 0.37579330801963811703;
            "LEFT_21_135": value  <= 0.66240137815475463867;
            "LEFT_21_136": value  <= 0.47957968711853027344;
            "LEFT_21_137": value  <= 0.49378821253776550293;
            "LEFT_21_138": value  <= 0.05389456078410150008;
            "LEFT_21_139": value  <= 0.51297742128372192383;
            "LEFT_21_140": value  <= 0.45283439755439758301;
            "LEFT_21_141": value  <= 0.53577268123626708984;
            "LEFT_21_142": value  <= 0.59161728620529174805;
            "LEFT_21_143": value  <= 0.52733850479125976562;
            "LEFT_21_144": value  <= 0.40465280413627630063;
            "LEFT_21_145": value  <= 0.74522358179092407227;
            "LEFT_21_146": value  <= 0.32954359054565429688;
            "LEFT_21_147": value  <= 0.48571440577507019043;
            "LEFT_21_148": value  <= 0.43127310276031488590;
            "LEFT_21_149": value  <= 0.51961702108383178711;
            "LEFT_21_150": value  <= 0.47357571125030517578;
            "LEFT_21_151": value  <= 0.58229267597198486328;
            "LEFT_21_152": value  <= 0.49991989135742187500;
            "LEFT_21_153": value  <= 0.47508931159973150082;
            "LEFT_21_154": value  <= 0.50697678327560424805;
            "LEFT_21_155": value  <= 0.48756939172744750977;
            "LEFT_21_156": value  <= 0.47507700324058532715;
            "LEFT_21_157": value  <= 0.53054618835449218750;
            "LEFT_21_158": value  <= 0.45184791088104248047;
            "LEFT_21_159": value  <= 0.41491198539733892270;
            "LEFT_21_160": value  <= 0.47178968787193298340;
            "LEFT_21_161": value  <= 0.21721640229225158691;
            "LEFT_21_162": value  <= 0.53373837471008300781;
            "LEFT_21_163": value  <= 0.46045941114425659180;
            "LEFT_21_164": value  <= 0.49458950757980352231;
            "LEFT_21_165": value  <= 0.70055091381072998047;
            "LEFT_21_166": value  <= 0.44662651419639587402;
            "LEFT_21_167": value  <= 0.47140988707542419434;
            "LEFT_21_168": value  <= 0.43315461277961730957;
            "LEFT_21_169": value  <= 0.26447001099586492368;
            "LEFT_21_170": value  <= 0.52083498239517211914;
            "LEFT_21_171": value  <= 0.63441252708435058594;
            "LEFT_21_172": value  <= 0.50504380464553833008;
            "LEFT_21_173": value  <= 0.49663180112838750668;
            "LEFT_21_174": value  <= 0.33002600073814392090;
            "LEFT_21_175": value  <= 0.49915981292724609375;
            "LEFT_21_176": value  <= 0.39117351174354547672;
            "LEFT_21_177": value  <= 0.56289112567901611328;
            "LEFT_21_178": value  <= 0.58535951375961303711;
            "LEFT_21_179": value  <= 0.42714700102806091309;
            "LEFT_21_180": value  <= 0.51431107521057128906;
            "LEFT_21_181": value  <= 0.60445022583007812500;
            "LEFT_21_182": value  <= 0.25831609964370727539;
            "LEFT_21_183": value  <= 0.48573741316795349121;
            "LEFT_21_184": value  <= 0.59368848800659179688;
            "LEFT_21_185": value  <= 0.31630149483680730649;
            "LEFT_21_186": value  <= 0.50612241029739379883;
            "LEFT_21_187": value  <= 0.47790178656578058414;
            "LEFT_21_188": value  <= 0.42978510260581970215;
            "LEFT_21_189": value  <= 0.54386717081069946289;
            "LEFT_21_190": value  <= 0.47268930077552800961;
            "LEFT_21_191": value  <= 0.42291730642318731137;
            "LEFT_21_192": value  <= 0.60988807678222656250;
            "LEFT_21_193": value  <= 0.56894367933273315430;
            "LEFT_21_194": value  <= 0.37622210383415222168;
            "LEFT_21_195": value  <= 0.46994051337242132016;
            "LEFT_21_196": value  <= 0.44652169942855840512;
            "LEFT_21_197": value  <= 0.54498052597045898438;
            "LEFT_21_198": value  <= 0.45640090107917791196;
            "LEFT_21_199": value  <= 0.57473778724670410156;
            "LEFT_21_200": value  <= 0.51661968231201171875;
            "LEFT_21_201": value  <= 0.50021117925643920898;
            "LEFT_21_202": value  <= 0.53945982456207275391;
            "LEFT_21_203": value  <= 0.51883268356323242188;
            "LEFT_21_204": value  <= 0.39046850800514221191;
            "LEFT_21_205": value  <= 0.48953229188919067383;
            "LEFT_21_206": value  <= 0.69752287864685058594;
            "LEFT_21_207": value  <= 0.52336359024047851562;
            "LEFT_21_208": value  <= 0.54193967580795288086;
            "LEFT_21_209": value  <= 0.48157641291618352719;
            "LEFT_21_210": value  <= 0.39802789688110351562;
            "LEFT_21_211": value  <= 0.54312318563461303711;
            "LEFT_21_212": value  <= 0.47382280230522161313;

            default: value <= -1;

        endcase

    end

endmodule 
