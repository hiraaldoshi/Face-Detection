module Width (

input int stage_num,
input int feature_num,
input int rectangle_num,
output real value

);

string name;
assign name = {"WIDTH_", $sformatf("%d", stage_num),
					"_", $sformatf("%d", feature_num), "_",
					$sformatf("%d", rectangle_num)};

always_comb
    begin

        case (name)

            "WIDTH_0_0_0": value  <=  14;
            "WIDTH_0_0_1": value  <=  14;
            "WIDTH_0_1_0": value  <=  18;
            "WIDTH_0_1_1": value  <=  6;
            "WIDTH_0_2_0": value  <=  15;
            "WIDTH_0_2_1": value  <=  15;
            "WIDTH_1_0_0": value  <=  2;
            "WIDTH_1_0_1": value  <=  2;
            "WIDTH_1_1_0": value  <=  6;
            "WIDTH_1_1_1": value  <=  2;
            "WIDTH_1_2_0": value  <=  12;
            "WIDTH_1_2_1": value  <=  12;
            "WIDTH_1_3_0": value  <=  10;
            "WIDTH_1_3_1": value  <=  10;
            "WIDTH_1_4_0": value  <=  14;
            "WIDTH_1_4_1": value  <=  14;
            "WIDTH_1_5_0": value  <=  6;
            "WIDTH_1_5_1": value  <=  3;
            "WIDTH_1_6_0": value  <=  5;
            "WIDTH_1_6_1": value  <=  5;
            "WIDTH_1_7_0": value  <=  18;
            "WIDTH_1_7_1": value  <=  6;
            "WIDTH_1_8_0": value  <=  17;
            "WIDTH_1_8_1": value  <=  17;
            "WIDTH_1_9_0": value  <=  4;
            "WIDTH_1_9_1": value  <=  4;
            "WIDTH_1_10_0": value  <=  2;
            "WIDTH_1_10_1": value  <=  2;
            "WIDTH_1_11_0": value  <=  6;
            "WIDTH_1_11_1": value  <=  3;
            "WIDTH_1_12_0": value  <=  4;
            "WIDTH_1_12_1": value  <=  2;
            "WIDTH_1_12_2": value  <=  2;
            "WIDTH_1_13_0": value  <=  18;
            "WIDTH_1_13_1": value  <=  6;
            "WIDTH_1_14_0": value  <=  10;
            "WIDTH_1_14_1": value  <=  10;
            "WIDTH_1_15_0": value  <=  5;
            "WIDTH_1_15_1": value  <=  5;
            "WIDTH_2_0_0": value  <=  10;
            "WIDTH_2_0_1": value  <=  10;
            "WIDTH_2_1_0": value  <=  2;
            "WIDTH_2_1_1": value  <=  2;
            "WIDTH_2_2_0": value  <=  4;
            "WIDTH_2_2_1": value  <=  4;
            "WIDTH_2_3_0": value  <=  12;
            "WIDTH_2_3_1": value  <=  4;
            "WIDTH_2_4_0": value  <=  10;
            "WIDTH_2_4_1": value  <=  10;
            "WIDTH_2_5_0": value  <=  6;
            "WIDTH_2_5_1": value  <=  6;
            "WIDTH_2_6_0": value  <=  1;
            "WIDTH_2_6_1": value  <=  1;
            "WIDTH_2_7_0": value  <=  20;
            "WIDTH_2_7_1": value  <=  20;
            "WIDTH_2_8_0": value  <=  6;
            "WIDTH_2_8_1": value  <=  2;
            "WIDTH_2_9_0": value  <=  6;
            "WIDTH_2_9_1": value  <=  2;
            "WIDTH_2_10_0": value  <=  6;
            "WIDTH_2_10_1": value  <=  2;
            "WIDTH_2_11_0": value  <=  6;
            "WIDTH_2_11_1": value  <=  2;
            "WIDTH_2_12_0": value  <=  18;
            "WIDTH_2_12_1": value  <=  9;
            "WIDTH_2_12_2": value  <=  9;
            "WIDTH_2_13_0": value  <=  10;
            "WIDTH_2_13_1": value  <=  5;
            "WIDTH_2_13_2": value  <=  5;
            "WIDTH_2_14_0": value  <=  4;
            "WIDTH_2_14_1": value  <=  2;
            "WIDTH_2_14_2": value  <=  2;
            "WIDTH_2_15_0": value  <=  14;
            "WIDTH_2_15_1": value  <=  7;
            "WIDTH_2_15_2": value  <=  7;
            "WIDTH_2_16_0": value  <=  6;
            "WIDTH_2_16_1": value  <=  2;
            "WIDTH_2_17_0": value  <=  20;
            "WIDTH_2_17_1": value  <=  20;
            "WIDTH_2_18_0": value  <=  4;
            "WIDTH_2_18_1": value  <=  4;
            "WIDTH_2_19_0": value  <=  2;
            "WIDTH_2_19_1": value  <=  2;
            "WIDTH_2_20_0": value  <=  9;
            "WIDTH_2_20_1": value  <=  9;
            "WIDTH_3_0_0": value  <=  3;
            "WIDTH_3_0_1": value  <=  3;
            "WIDTH_3_1_0": value  <=  2;
            "WIDTH_3_1_1": value  <=  2;
            "WIDTH_3_2_0": value  <=  13;
            "WIDTH_3_2_1": value  <=  13;
            "WIDTH_3_3_0": value  <=  8;
            "WIDTH_3_3_1": value  <=  4;
            "WIDTH_3_4_0": value  <=  4;
            "WIDTH_3_4_1": value  <=  4;
            "WIDTH_3_5_0": value  <=  8;
            "WIDTH_3_5_1": value  <=  4;
            "WIDTH_3_5_2": value  <=  4;
            "WIDTH_3_6_0": value  <=  6;
            "WIDTH_3_6_1": value  <=  2;
            "WIDTH_3_7_0": value  <=  6;
            "WIDTH_3_7_1": value  <=  2;
            "WIDTH_3_8_0": value  <=  9;
            "WIDTH_3_8_1": value  <=  3;
            "WIDTH_3_9_0": value  <=  10;
            "WIDTH_3_9_1": value  <=  5;
            "WIDTH_3_9_2": value  <=  5;
            "WIDTH_3_10_0": value  <=  6;
            "WIDTH_3_10_1": value  <=  3;
            "WIDTH_3_11_0": value  <=  15;
            "WIDTH_3_11_1": value  <=  15;
            "WIDTH_3_12_0": value  <=  8;
            "WIDTH_3_12_1": value  <=  8;
            "WIDTH_3_13_0": value  <=  12;
            "WIDTH_3_13_1": value  <=  6;
            "WIDTH_3_13_2": value  <=  6;
            "WIDTH_3_14_0": value  <=  4;
            "WIDTH_3_14_1": value  <=  2;
            "WIDTH_3_15_0": value  <=  1;
            "WIDTH_3_15_1": value  <=  1;
            "WIDTH_3_16_0": value  <=  2;
            "WIDTH_3_16_1": value  <=  2;
            "WIDTH_3_17_0": value  <=  1;
            "WIDTH_3_17_1": value  <=  1;
            "WIDTH_3_18_0": value  <=  6;
            "WIDTH_3_18_1": value  <=  3;
            "WIDTH_3_18_2": value  <=  3;
            "WIDTH_3_19_0": value  <=  8;
            "WIDTH_3_19_1": value  <=  8;
            "WIDTH_3_20_0": value  <=  1;
            "WIDTH_3_20_1": value  <=  1;
            "WIDTH_3_21_0": value  <=  12;
            "WIDTH_3_21_1": value  <=  12;
            "WIDTH_3_22_0": value  <=  2;
            "WIDTH_3_22_1": value  <=  2;
            "WIDTH_3_23_0": value  <=  6;
            "WIDTH_3_23_1": value  <=  6;
            "WIDTH_3_24_0": value  <=  4;
            "WIDTH_3_24_1": value  <=  4;
            "WIDTH_3_25_0": value  <=  12;
            "WIDTH_3_25_1": value  <=  4;
            "WIDTH_3_26_0": value  <=  1;
            "WIDTH_3_26_1": value  <=  1;
            "WIDTH_3_27_0": value  <=  3;
            "WIDTH_3_27_1": value  <=  1;
            "WIDTH_3_28_0": value  <=  2;
            "WIDTH_3_28_1": value  <=  2;
            "WIDTH_3_29_0": value  <=  6;
            "WIDTH_3_29_1": value  <=  2;
            "WIDTH_3_30_0": value  <=  3;
            "WIDTH_3_30_1": value  <=  1;
            "WIDTH_3_31_0": value  <=  3;
            "WIDTH_3_31_1": value  <=  1;
            "WIDTH_3_32_0": value  <=  3;
            "WIDTH_3_32_1": value  <=  3;
            "WIDTH_3_33_0": value  <=  6;
            "WIDTH_3_33_1": value  <=  2;
            "WIDTH_3_34_0": value  <=  14;
            "WIDTH_3_34_1": value  <=  14;
            "WIDTH_3_35_0": value  <=  18;
            "WIDTH_3_35_1": value  <=  9;
            "WIDTH_3_35_2": value  <=  9;
            "WIDTH_3_36_0": value  <=  3;
            "WIDTH_3_36_1": value  <=  3;
            "WIDTH_3_37_0": value  <=  6;
            "WIDTH_3_37_1": value  <=  2;
            "WIDTH_3_38_0": value  <=  3;
            "WIDTH_3_38_1": value  <=  1;
            "WIDTH_4_0_0": value  <=  18;
            "WIDTH_4_0_1": value  <=  18;
            "WIDTH_4_1_0": value  <=  2;
            "WIDTH_4_1_1": value  <=  2;
            "WIDTH_4_2_0": value  <=  19;
            "WIDTH_4_2_1": value  <=  19;
            "WIDTH_4_3_0": value  <=  6;
            "WIDTH_4_3_1": value  <=  2;
            "WIDTH_4_4_0": value  <=  6;
            "WIDTH_4_4_1": value  <=  2;
            "WIDTH_4_5_0": value  <=  6;
            "WIDTH_4_5_1": value  <=  2;
            "WIDTH_4_6_0": value  <=  4;
            "WIDTH_4_6_1": value  <=  4;
            "WIDTH_4_7_0": value  <=  6;
            "WIDTH_4_7_1": value  <=  2;
            "WIDTH_4_8_0": value  <=  12;
            "WIDTH_4_8_1": value  <=  12;
            "WIDTH_4_9_0": value  <=  2;
            "WIDTH_4_9_1": value  <=  2;
            "WIDTH_4_10_0": value  <=  2;
            "WIDTH_4_10_1": value  <=  1;
            "WIDTH_4_11_0": value  <=  3;
            "WIDTH_4_11_1": value  <=  1;
            "WIDTH_4_12_0": value  <=  4;
            "WIDTH_4_12_1": value  <=  2;
            "WIDTH_4_13_0": value  <=  4;
            "WIDTH_4_13_1": value  <=  2;
            "WIDTH_4_13_2": value  <=  2;
            "WIDTH_4_14_0": value  <=  1;
            "WIDTH_4_14_1": value  <=  1;
            "WIDTH_4_15_0": value  <=  1;
            "WIDTH_4_15_1": value  <=  1;
            "WIDTH_4_16_0": value  <=  6;
            "WIDTH_4_16_1": value  <=  3;
            "WIDTH_4_17_0": value  <=  3;
            "WIDTH_4_17_1": value  <=  1;
            "WIDTH_4_18_0": value  <=  3;
            "WIDTH_4_18_1": value  <=  1;
            "WIDTH_4_19_0": value  <=  12;
            "WIDTH_4_19_1": value  <=  12;
            "WIDTH_4_20_0": value  <=  2;
            "WIDTH_4_20_1": value  <=  2;
            "WIDTH_4_21_0": value  <=  2;
            "WIDTH_4_21_1": value  <=  2;
            "WIDTH_4_22_0": value  <=  3;
            "WIDTH_4_22_1": value  <=  1;
            "WIDTH_4_23_0": value  <=  6;
            "WIDTH_4_23_1": value  <=  2;
            "WIDTH_4_24_0": value  <=  9;
            "WIDTH_4_24_1": value  <=  9;
            "WIDTH_4_25_0": value  <=  6;
            "WIDTH_4_25_1": value  <=  2;
            "WIDTH_4_26_0": value  <=  18;
            "WIDTH_4_26_1": value  <=  6;
            "WIDTH_4_27_0": value  <=  4;
            "WIDTH_4_27_1": value  <=  2;
            "WIDTH_4_27_2": value  <=  2;
            "WIDTH_4_28_0": value  <=  1;
            "WIDTH_4_28_1": value  <=  1;
            "WIDTH_4_29_0": value  <=  5;
            "WIDTH_4_29_1": value  <=  5;
            "WIDTH_4_30_0": value  <=  10;
            "WIDTH_4_30_1": value  <=  5;
            "WIDTH_4_30_2": value  <=  5;
            "WIDTH_4_31_0": value  <=  9;
            "WIDTH_4_31_1": value  <=  9;
            "WIDTH_4_32_0": value  <=  12;
            "WIDTH_4_32_1": value  <=  6;
            "WIDTH_4_32_2": value  <=  6;
            "WIDTH_5_0_0": value  <=  12;
            "WIDTH_5_0_1": value  <=  4;
            "WIDTH_5_1_0": value  <=  6;
            "WIDTH_5_1_1": value  <=  6;
            "WIDTH_5_2_0": value  <=  11;
            "WIDTH_5_2_1": value  <=  11;
            "WIDTH_5_3_0": value  <=  16;
            "WIDTH_5_3_1": value  <=  16;
            "WIDTH_5_4_0": value  <=  16;
            "WIDTH_5_4_1": value  <=  16;
            "WIDTH_5_5_0": value  <=  6;
            "WIDTH_5_5_1": value  <=  2;
            "WIDTH_5_6_0": value  <=  6;
            "WIDTH_5_6_1": value  <=  3;
            "WIDTH_5_6_2": value  <=  3;
            "WIDTH_5_7_0": value  <=  8;
            "WIDTH_5_7_1": value  <=  8;
            "WIDTH_5_8_0": value  <=  8;
            "WIDTH_5_8_1": value  <=  4;
            "WIDTH_5_8_2": value  <=  4;
            "WIDTH_5_9_0": value  <=  2;
            "WIDTH_5_9_1": value  <=  2;
            "WIDTH_5_10_0": value  <=  7;
            "WIDTH_5_10_1": value  <=  7;
            "WIDTH_5_11_0": value  <=  4;
            "WIDTH_5_11_1": value  <=  2;
            "WIDTH_5_12_0": value  <=  14;
            "WIDTH_5_12_1": value  <=  7;
            "WIDTH_5_12_2": value  <=  7;
            "WIDTH_5_13_0": value  <=  10;
            "WIDTH_5_13_1": value  <=  10;
            "WIDTH_5_14_0": value  <=  8;
            "WIDTH_5_14_1": value  <=  4;
            "WIDTH_5_14_2": value  <=  4;
            "WIDTH_5_15_0": value  <=  3;
            "WIDTH_5_15_1": value  <=  3;
            "WIDTH_5_16_0": value  <=  4;
            "WIDTH_5_16_1": value  <=  2;
            "WIDTH_5_17_0": value  <=  2;
            "WIDTH_5_17_1": value  <=  2;
            "WIDTH_5_18_0": value  <=  5;
            "WIDTH_5_18_1": value  <=  5;
            "WIDTH_5_19_0": value  <=  18;
            "WIDTH_5_19_1": value  <=  9;
            "WIDTH_5_19_2": value  <=  9;
            "WIDTH_5_20_0": value  <=  1;
            "WIDTH_5_20_1": value  <=  1;
            "WIDTH_5_21_0": value  <=  1;
            "WIDTH_5_21_1": value  <=  1;
            "WIDTH_5_22_0": value  <=  6;
            "WIDTH_5_22_1": value  <=  2;
            "WIDTH_5_23_0": value  <=  1;
            "WIDTH_5_23_1": value  <=  1;
            "WIDTH_5_24_0": value  <=  2;
            "WIDTH_5_24_1": value  <=  2;
            "WIDTH_5_25_0": value  <=  8;
            "WIDTH_5_25_1": value  <=  4;
            "WIDTH_5_25_2": value  <=  4;
            "WIDTH_5_26_0": value  <=  6;
            "WIDTH_5_26_1": value  <=  2;
            "WIDTH_5_27_0": value  <=  9;
            "WIDTH_5_27_1": value  <=  9;
            "WIDTH_5_28_0": value  <=  6;
            "WIDTH_5_28_1": value  <=  2;
            "WIDTH_5_29_0": value  <=  2;
            "WIDTH_5_29_1": value  <=  2;
            "WIDTH_5_30_0": value  <=  5;
            "WIDTH_5_30_1": value  <=  5;
            "WIDTH_5_31_0": value  <=  3;
            "WIDTH_5_31_1": value  <=  3;
            "WIDTH_5_32_0": value  <=  8;
            "WIDTH_5_32_1": value  <=  8;
            "WIDTH_5_33_0": value  <=  3;
            "WIDTH_5_33_1": value  <=  3;
            "WIDTH_5_34_0": value  <=  3;
            "WIDTH_5_34_1": value  <=  3;
            "WIDTH_5_35_0": value  <=  12;
            "WIDTH_5_35_1": value  <=  6;
            "WIDTH_5_35_2": value  <=  6;
            "WIDTH_5_36_0": value  <=  2;
            "WIDTH_5_36_1": value  <=  1;
            "WIDTH_5_37_0": value  <=  5;
            "WIDTH_5_37_1": value  <=  5;
            "WIDTH_5_38_0": value  <=  3;
            "WIDTH_5_38_1": value  <=  1;
            "WIDTH_5_39_0": value  <=  2;
            "WIDTH_5_39_1": value  <=  2;
            "WIDTH_5_40_0": value  <=  3;
            "WIDTH_5_40_1": value  <=  1;
            "WIDTH_5_41_0": value  <=  3;
            "WIDTH_5_41_1": value  <=  1;
            "WIDTH_5_42_0": value  <=  6;
            "WIDTH_5_42_1": value  <=  2;
            "WIDTH_5_43_0": value  <=  10;
            "WIDTH_5_43_1": value  <=  10;
            "WIDTH_6_0_0": value  <=  6;
            "WIDTH_6_0_1": value  <=  6;
            "WIDTH_6_1_0": value  <=  9;
            "WIDTH_6_1_1": value  <=  3;
            "WIDTH_6_2_0": value  <=  16;
            "WIDTH_6_2_1": value  <=  16;
            "WIDTH_6_3_0": value  <=  2;
            "WIDTH_6_3_1": value  <=  2;
            "WIDTH_6_4_0": value  <=  6;
            "WIDTH_6_4_1": value  <=  6;
            "WIDTH_6_5_0": value  <=  6;
            "WIDTH_6_5_1": value  <=  6;
            "WIDTH_6_6_0": value  <=  7;
            "WIDTH_6_6_1": value  <=  7;
            "WIDTH_6_7_0": value  <=  3;
            "WIDTH_6_7_1": value  <=  3;
            "WIDTH_6_8_0": value  <=  15;
            "WIDTH_6_8_1": value  <=  5;
            "WIDTH_6_9_0": value  <=  3;
            "WIDTH_6_9_1": value  <=  3;
            "WIDTH_6_10_0": value  <=  4;
            "WIDTH_6_10_1": value  <=  4;
            "WIDTH_6_11_0": value  <=  6;
            "WIDTH_6_11_1": value  <=  2;
            "WIDTH_6_12_0": value  <=  8;
            "WIDTH_6_12_1": value  <=  4;
            "WIDTH_6_12_2": value  <=  4;
            "WIDTH_6_13_0": value  <=  12;
            "WIDTH_6_13_1": value  <=  6;
            "WIDTH_6_13_2": value  <=  6;
            "WIDTH_6_14_0": value  <=  6;
            "WIDTH_6_14_1": value  <=  2;
            "WIDTH_6_15_0": value  <=  2;
            "WIDTH_6_15_1": value  <=  1;
            "WIDTH_6_16_0": value  <=  2;
            "WIDTH_6_16_1": value  <=  1;
            "WIDTH_6_17_0": value  <=  2;
            "WIDTH_6_17_1": value  <=  2;
            "WIDTH_6_18_0": value  <=  6;
            "WIDTH_6_18_1": value  <=  3;
            "WIDTH_6_19_0": value  <=  2;
            "WIDTH_6_19_1": value  <=  2;
            "WIDTH_6_20_0": value  <=  12;
            "WIDTH_6_20_1": value  <=  12;
            "WIDTH_6_21_0": value  <=  5;
            "WIDTH_6_21_1": value  <=  5;
            "WIDTH_6_22_0": value  <=  3;
            "WIDTH_6_22_1": value  <=  3;
            "WIDTH_6_23_0": value  <=  3;
            "WIDTH_6_23_1": value  <=  1;
            "WIDTH_6_24_0": value  <=  6;
            "WIDTH_6_24_1": value  <=  3;
            "WIDTH_6_25_0": value  <=  1;
            "WIDTH_6_25_1": value  <=  1;
            "WIDTH_6_26_0": value  <=  4;
            "WIDTH_6_26_1": value  <=  2;
            "WIDTH_6_26_2": value  <=  2;
            "WIDTH_6_27_0": value  <=  4;
            "WIDTH_6_27_1": value  <=  4;
            "WIDTH_6_28_0": value  <=  4;
            "WIDTH_6_28_1": value  <=  4;
            "WIDTH_6_29_0": value  <=  3;
            "WIDTH_6_29_1": value  <=  3;
            "WIDTH_6_30_0": value  <=  4;
            "WIDTH_6_30_1": value  <=  4;
            "WIDTH_6_31_0": value  <=  11;
            "WIDTH_6_31_1": value  <=  11;
            "WIDTH_6_32_0": value  <=  3;
            "WIDTH_6_32_1": value  <=  1;
            "WIDTH_6_33_0": value  <=  6;
            "WIDTH_6_33_1": value  <=  2;
            "WIDTH_6_34_0": value  <=  3;
            "WIDTH_6_34_1": value  <=  3;
            "WIDTH_6_35_0": value  <=  20;
            "WIDTH_6_35_1": value  <=  10;
            "WIDTH_6_35_2": value  <=  10;
            "WIDTH_6_36_0": value  <=  3;
            "WIDTH_6_36_1": value  <=  1;
            "WIDTH_6_37_0": value  <=  1;
            "WIDTH_6_37_1": value  <=  1;
            "WIDTH_6_38_0": value  <=  4;
            "WIDTH_6_38_1": value  <=  4;
            "WIDTH_6_39_0": value  <=  4;
            "WIDTH_6_39_1": value  <=  4;
            "WIDTH_6_40_0": value  <=  6;
            "WIDTH_6_40_1": value  <=  2;
            "WIDTH_6_41_0": value  <=  3;
            "WIDTH_6_41_1": value  <=  1;
            "WIDTH_6_42_0": value  <=  2;
            "WIDTH_6_42_1": value  <=  1;
            "WIDTH_6_43_0": value  <=  14;
            "WIDTH_6_43_1": value  <=  7;
            "WIDTH_6_43_2": value  <=  7;
            "WIDTH_6_44_0": value  <=  3;
            "WIDTH_6_44_1": value  <=  3;
            "WIDTH_6_45_0": value  <=  3;
            "WIDTH_6_45_1": value  <=  3;
            "WIDTH_6_46_0": value  <=  3;
            "WIDTH_6_46_1": value  <=  3;
            "WIDTH_6_47_0": value  <=  12;
            "WIDTH_6_47_1": value  <=  6;
            "WIDTH_6_47_2": value  <=  6;
            "WIDTH_6_48_0": value  <=  1;
            "WIDTH_6_48_1": value  <=  1;
            "WIDTH_6_49_0": value  <=  2;
            "WIDTH_6_49_1": value  <=  2;
            "WIDTH_7_0_0": value  <=  6;
            "WIDTH_7_0_1": value  <=  2;
            "WIDTH_7_1_0": value  <=  6;
            "WIDTH_7_1_1": value  <=  3;
            "WIDTH_7_1_2": value  <=  3;
            "WIDTH_7_2_0": value  <=  10;
            "WIDTH_7_2_1": value  <=  10;
            "WIDTH_7_3_0": value  <=  8;
            "WIDTH_7_3_1": value  <=  4;
            "WIDTH_7_3_2": value  <=  4;
            "WIDTH_7_4_0": value  <=  7;
            "WIDTH_7_4_1": value  <=  7;
            "WIDTH_7_5_0": value  <=  6;
            "WIDTH_7_5_1": value  <=  3;
            "WIDTH_7_5_2": value  <=  3;
            "WIDTH_7_6_0": value  <=  6;
            "WIDTH_7_6_1": value  <=  3;
            "WIDTH_7_6_2": value  <=  3;
            "WIDTH_7_7_0": value  <=  18;
            "WIDTH_7_7_1": value  <=  6;
            "WIDTH_7_8_0": value  <=  8;
            "WIDTH_7_8_1": value  <=  4;
            "WIDTH_7_8_2": value  <=  4;
            "WIDTH_7_9_0": value  <=  2;
            "WIDTH_7_9_1": value  <=  2;
            "WIDTH_7_10_0": value  <=  2;
            "WIDTH_7_10_1": value  <=  2;
            "WIDTH_7_11_0": value  <=  2;
            "WIDTH_7_11_1": value  <=  2;
            "WIDTH_7_12_0": value  <=  2;
            "WIDTH_7_12_1": value  <=  2;
            "WIDTH_7_13_0": value  <=  18;
            "WIDTH_7_13_1": value  <=  18;
            "WIDTH_7_14_0": value  <=  6;
            "WIDTH_7_14_1": value  <=  3;
            "WIDTH_7_15_0": value  <=  6;
            "WIDTH_7_15_1": value  <=  6;
            "WIDTH_7_16_0": value  <=  13;
            "WIDTH_7_16_1": value  <=  13;
            "WIDTH_7_17_0": value  <=  2;
            "WIDTH_7_17_1": value  <=  2;
            "WIDTH_7_18_0": value  <=  16;
            "WIDTH_7_18_1": value  <=  8;
            "WIDTH_7_18_2": value  <=  8;
            "WIDTH_7_19_0": value  <=  6;
            "WIDTH_7_19_1": value  <=  3;
            "WIDTH_7_19_2": value  <=  3;
            "WIDTH_7_20_0": value  <=  3;
            "WIDTH_7_20_1": value  <=  3;
            "WIDTH_7_21_0": value  <=  1;
            "WIDTH_7_21_1": value  <=  1;
            "WIDTH_7_22_0": value  <=  4;
            "WIDTH_7_22_1": value  <=  2;
            "WIDTH_7_23_0": value  <=  15;
            "WIDTH_7_23_1": value  <=  5;
            "WIDTH_7_24_0": value  <=  5;
            "WIDTH_7_24_1": value  <=  5;
            "WIDTH_7_25_0": value  <=  17;
            "WIDTH_7_25_1": value  <=  17;
            "WIDTH_7_26_0": value  <=  8;
            "WIDTH_7_26_1": value  <=  4;
            "WIDTH_7_27_0": value  <=  3;
            "WIDTH_7_27_1": value  <=  1;
            "WIDTH_7_28_0": value  <=  3;
            "WIDTH_7_28_1": value  <=  1;
            "WIDTH_7_29_0": value  <=  4;
            "WIDTH_7_29_1": value  <=  4;
            "WIDTH_7_30_0": value  <=  4;
            "WIDTH_7_30_1": value  <=  4;
            "WIDTH_7_31_0": value  <=  6;
            "WIDTH_7_31_1": value  <=  3;
            "WIDTH_7_32_0": value  <=  4;
            "WIDTH_7_32_1": value  <=  4;
            "WIDTH_7_33_0": value  <=  12;
            "WIDTH_7_33_1": value  <=  6;
            "WIDTH_7_33_2": value  <=  6;
            "WIDTH_7_34_0": value  <=  4;
            "WIDTH_7_34_1": value  <=  4;
            "WIDTH_7_35_0": value  <=  3;
            "WIDTH_7_35_1": value  <=  3;
            "WIDTH_7_36_0": value  <=  3;
            "WIDTH_7_36_1": value  <=  1;
            "WIDTH_7_37_0": value  <=  3;
            "WIDTH_7_37_1": value  <=  1;
            "WIDTH_7_38_0": value  <=  4;
            "WIDTH_7_38_1": value  <=  2;
            "WIDTH_7_39_0": value  <=  6;
            "WIDTH_7_39_1": value  <=  3;
            "WIDTH_7_40_0": value  <=  3;
            "WIDTH_7_40_1": value  <=  3;
            "WIDTH_7_41_0": value  <=  6;
            "WIDTH_7_41_1": value  <=  3;
            "WIDTH_7_42_0": value  <=  10;
            "WIDTH_7_42_1": value  <=  5;
            "WIDTH_7_42_2": value  <=  5;
            "WIDTH_7_43_0": value  <=  6;
            "WIDTH_7_43_1": value  <=  3;
            "WIDTH_7_44_0": value  <=  6;
            "WIDTH_7_44_1": value  <=  3;
            "WIDTH_7_45_0": value  <=  4;
            "WIDTH_7_45_1": value  <=  2;
            "WIDTH_7_46_0": value  <=  2;
            "WIDTH_7_46_1": value  <=  1;
            "WIDTH_7_47_0": value  <=  4;
            "WIDTH_7_47_1": value  <=  2;
            "WIDTH_7_47_2": value  <=  2;
            "WIDTH_7_48_0": value  <=  2;
            "WIDTH_7_48_1": value  <=  1;
            "WIDTH_7_49_0": value  <=  12;
            "WIDTH_7_49_1": value  <=  4;
            "WIDTH_7_50_0": value  <=  3;
            "WIDTH_7_50_1": value  <=  1;
            "WIDTH_8_0_0": value  <=  8;
            "WIDTH_8_0_1": value  <=  8;
            "WIDTH_8_1_0": value  <=  2;
            "WIDTH_8_1_1": value  <=  2;
            "WIDTH_8_2_0": value  <=  6;
            "WIDTH_8_2_1": value  <=  6;
            "WIDTH_8_3_0": value  <=  8;
            "WIDTH_8_3_1": value  <=  4;
            "WIDTH_8_4_0": value  <=  18;
            "WIDTH_8_4_1": value  <=  18;
            "WIDTH_8_5_0": value  <=  4;
            "WIDTH_8_5_1": value  <=  4;
            "WIDTH_8_6_0": value  <=  8;
            "WIDTH_8_6_1": value  <=  4;
            "WIDTH_8_7_0": value  <=  3;
            "WIDTH_8_7_1": value  <=  3;
            "WIDTH_8_8_0": value  <=  6;
            "WIDTH_8_8_1": value  <=  2;
            "WIDTH_8_9_0": value  <=  3;
            "WIDTH_8_9_1": value  <=  1;
            "WIDTH_8_10_0": value  <=  5;
            "WIDTH_8_10_1": value  <=  5;
            "WIDTH_8_11_0": value  <=  7;
            "WIDTH_8_11_1": value  <=  7;
            "WIDTH_8_12_0": value  <=  7;
            "WIDTH_8_12_1": value  <=  7;
            "WIDTH_8_13_0": value  <=  2;
            "WIDTH_8_13_1": value  <=  2;
            "WIDTH_8_14_0": value  <=  3;
            "WIDTH_8_14_1": value  <=  3;
            "WIDTH_8_15_0": value  <=  3;
            "WIDTH_8_15_1": value  <=  1;
            "WIDTH_8_16_0": value  <=  4;
            "WIDTH_8_16_1": value  <=  2;
            "WIDTH_8_17_0": value  <=  6;
            "WIDTH_8_17_1": value  <=  2;
            "WIDTH_8_18_0": value  <=  3;
            "WIDTH_8_18_1": value  <=  3;
            "WIDTH_8_19_0": value  <=  4;
            "WIDTH_8_19_1": value  <=  4;
            "WIDTH_8_20_0": value  <=  4;
            "WIDTH_8_20_1": value  <=  4;
            "WIDTH_8_21_0": value  <=  18;
            "WIDTH_8_21_1": value  <=  18;
            "WIDTH_8_22_0": value  <=  3;
            "WIDTH_8_22_1": value  <=  1;
            "WIDTH_8_23_0": value  <=  6;
            "WIDTH_8_23_1": value  <=  3;
            "WIDTH_8_23_2": value  <=  3;
            "WIDTH_8_24_0": value  <=  3;
            "WIDTH_8_24_1": value  <=  3;
            "WIDTH_8_25_0": value  <=  20;
            "WIDTH_8_25_1": value  <=  10;
            "WIDTH_8_25_2": value  <=  10;
            "WIDTH_8_26_0": value  <=  6;
            "WIDTH_8_26_1": value  <=  2;
            "WIDTH_8_27_0": value  <=  2;
            "WIDTH_8_27_1": value  <=  2;
            "WIDTH_8_28_0": value  <=  6;
            "WIDTH_8_28_1": value  <=  3;
            "WIDTH_8_28_2": value  <=  3;
            "WIDTH_8_29_0": value  <=  20;
            "WIDTH_8_29_1": value  <=  10;
            "WIDTH_8_29_2": value  <=  10;
            "WIDTH_8_30_0": value  <=  5;
            "WIDTH_8_30_1": value  <=  5;
            "WIDTH_8_31_0": value  <=  6;
            "WIDTH_8_31_1": value  <=  3;
            "WIDTH_8_31_2": value  <=  3;
            "WIDTH_8_32_0": value  <=  2;
            "WIDTH_8_32_1": value  <=  2;
            "WIDTH_8_33_0": value  <=  1;
            "WIDTH_8_33_1": value  <=  1;
            "WIDTH_8_34_0": value  <=  1;
            "WIDTH_8_34_1": value  <=  1;
            "WIDTH_8_35_0": value  <=  14;
            "WIDTH_8_35_1": value  <=  7;
            "WIDTH_8_35_2": value  <=  7;
            "WIDTH_8_36_0": value  <=  3;
            "WIDTH_8_36_1": value  <=  3;
            "WIDTH_8_37_0": value  <=  3;
            "WIDTH_8_37_1": value  <=  1;
            "WIDTH_8_38_0": value  <=  8;
            "WIDTH_8_38_1": value  <=  8;
            "WIDTH_8_39_0": value  <=  3;
            "WIDTH_8_39_1": value  <=  1;
            "WIDTH_8_40_0": value  <=  4;
            "WIDTH_8_40_1": value  <=  2;
            "WIDTH_8_40_2": value  <=  2;
            "WIDTH_8_41_0": value  <=  10;
            "WIDTH_8_41_1": value  <=  5;
            "WIDTH_8_42_0": value  <=  3;
            "WIDTH_8_42_1": value  <=  1;
            "WIDTH_8_43_0": value  <=  2;
            "WIDTH_8_43_1": value  <=  2;
            "WIDTH_8_44_0": value  <=  3;
            "WIDTH_8_44_1": value  <=  1;
            "WIDTH_8_45_0": value  <=  1;
            "WIDTH_8_45_1": value  <=  1;
            "WIDTH_8_46_0": value  <=  12;
            "WIDTH_8_46_1": value  <=  6;
            "WIDTH_8_46_2": value  <=  6;
            "WIDTH_8_47_0": value  <=  7;
            "WIDTH_8_47_1": value  <=  7;
            "WIDTH_8_48_0": value  <=  2;
            "WIDTH_8_48_1": value  <=  2;
            "WIDTH_8_49_0": value  <=  14;
            "WIDTH_8_49_1": value  <=  7;
            "WIDTH_8_49_2": value  <=  7;
            "WIDTH_8_50_0": value  <=  3;
            "WIDTH_8_50_1": value  <=  1;
            "WIDTH_8_51_0": value  <=  6;
            "WIDTH_8_51_1": value  <=  2;
            "WIDTH_8_52_0": value  <=  6;
            "WIDTH_8_52_1": value  <=  3;
            "WIDTH_8_53_0": value  <=  6;
            "WIDTH_8_53_1": value  <=  6;
            "WIDTH_8_54_0": value  <=  18;
            "WIDTH_8_54_1": value  <=  6;
            "WIDTH_8_55_0": value  <=  3;
            "WIDTH_8_55_1": value  <=  3;
            "WIDTH_9_0_0": value  <=  7;
            "WIDTH_9_0_1": value  <=  7;
            "WIDTH_9_1_0": value  <=  12;
            "WIDTH_9_1_1": value  <=  4;
            "WIDTH_9_2_0": value  <=  17;
            "WIDTH_9_2_1": value  <=  17;
            "WIDTH_9_3_0": value  <=  15;
            "WIDTH_9_3_1": value  <=  15;
            "WIDTH_9_4_0": value  <=  6;
            "WIDTH_9_4_1": value  <=  6;
            "WIDTH_9_5_0": value  <=  4;
            "WIDTH_9_5_1": value  <=  2;
            "WIDTH_9_6_0": value  <=  3;
            "WIDTH_9_6_1": value  <=  3;
            "WIDTH_9_7_0": value  <=  7;
            "WIDTH_9_7_1": value  <=  7;
            "WIDTH_9_8_0": value  <=  4;
            "WIDTH_9_8_1": value  <=  4;
            "WIDTH_9_9_0": value  <=  20;
            "WIDTH_9_9_1": value  <=  10;
            "WIDTH_9_9_2": value  <=  10;
            "WIDTH_9_10_0": value  <=  6;
            "WIDTH_9_10_1": value  <=  3;
            "WIDTH_9_10_2": value  <=  3;
            "WIDTH_9_11_0": value  <=  3;
            "WIDTH_9_11_1": value  <=  3;
            "WIDTH_9_12_0": value  <=  3;
            "WIDTH_9_12_1": value  <=  3;
            "WIDTH_9_13_0": value  <=  6;
            "WIDTH_9_13_1": value  <=  2;
            "WIDTH_9_14_0": value  <=  6;
            "WIDTH_9_14_1": value  <=  6;
            "WIDTH_9_15_0": value  <=  20;
            "WIDTH_9_15_1": value  <=  20;
            "WIDTH_9_16_0": value  <=  4;
            "WIDTH_9_16_1": value  <=  2;
            "WIDTH_9_16_2": value  <=  2;
            "WIDTH_9_17_0": value  <=  8;
            "WIDTH_9_17_1": value  <=  4;
            "WIDTH_9_17_2": value  <=  4;
            "WIDTH_9_18_0": value  <=  15;
            "WIDTH_9_18_1": value  <=  15;
            "WIDTH_9_19_0": value  <=  2;
            "WIDTH_9_19_1": value  <=  2;
            "WIDTH_9_20_0": value  <=  1;
            "WIDTH_9_20_1": value  <=  1;
            "WIDTH_9_21_0": value  <=  2;
            "WIDTH_9_21_1": value  <=  2;
            "WIDTH_9_22_0": value  <=  3;
            "WIDTH_9_22_1": value  <=  1;
            "WIDTH_9_23_0": value  <=  3;
            "WIDTH_9_23_1": value  <=  3;
            "WIDTH_9_24_0": value  <=  3;
            "WIDTH_9_24_1": value  <=  1;
            "WIDTH_9_25_0": value  <=  5;
            "WIDTH_9_25_1": value  <=  5;
            "WIDTH_9_26_0": value  <=  5;
            "WIDTH_9_26_1": value  <=  5;
            "WIDTH_9_27_0": value  <=  1;
            "WIDTH_9_27_1": value  <=  1;
            "WIDTH_9_28_0": value  <=  4;
            "WIDTH_9_28_1": value  <=  4;
            "WIDTH_9_29_0": value  <=  3;
            "WIDTH_9_29_1": value  <=  3;
            "WIDTH_9_30_0": value  <=  3;
            "WIDTH_9_30_1": value  <=  3;
            "WIDTH_9_31_0": value  <=  6;
            "WIDTH_9_31_1": value  <=  6;
            "WIDTH_9_32_0": value  <=  5;
            "WIDTH_9_32_1": value  <=  5;
            "WIDTH_9_33_0": value  <=  6;
            "WIDTH_9_33_1": value  <=  2;
            "WIDTH_9_34_0": value  <=  6;
            "WIDTH_9_34_1": value  <=  2;
            "WIDTH_9_35_0": value  <=  4;
            "WIDTH_9_35_1": value  <=  4;
            "WIDTH_9_36_0": value  <=  3;
            "WIDTH_9_36_1": value  <=  3;
            "WIDTH_9_37_0": value  <=  8;
            "WIDTH_9_37_1": value  <=  8;
            "WIDTH_9_38_0": value  <=  5;
            "WIDTH_9_38_1": value  <=  5;
            "WIDTH_9_39_0": value  <=  4;
            "WIDTH_9_39_1": value  <=  2;
            "WIDTH_9_40_0": value  <=  3;
            "WIDTH_9_40_1": value  <=  3;
            "WIDTH_9_41_0": value  <=  1;
            "WIDTH_9_41_1": value  <=  1;
            "WIDTH_9_42_0": value  <=  4;
            "WIDTH_9_42_1": value  <=  2;
            "WIDTH_9_43_0": value  <=  4;
            "WIDTH_9_43_1": value  <=  2;
            "WIDTH_9_44_0": value  <=  4;
            "WIDTH_9_44_1": value  <=  2;
            "WIDTH_9_45_0": value  <=  15;
            "WIDTH_9_45_1": value  <=  5;
            "WIDTH_9_46_0": value  <=  6;
            "WIDTH_9_46_1": value  <=  3;
            "WIDTH_9_47_0": value  <=  3;
            "WIDTH_9_47_1": value  <=  1;
            "WIDTH_9_48_0": value  <=  3;
            "WIDTH_9_48_1": value  <=  3;
            "WIDTH_9_49_0": value  <=  5;
            "WIDTH_9_49_1": value  <=  5;
            "WIDTH_9_50_0": value  <=  4;
            "WIDTH_9_50_1": value  <=  4;
            "WIDTH_9_51_0": value  <=  3;
            "WIDTH_9_51_1": value  <=  1;
            "WIDTH_9_52_0": value  <=  14;
            "WIDTH_9_52_1": value  <=  7;
            "WIDTH_9_52_2": value  <=  7;
            "WIDTH_9_53_0": value  <=  16;
            "WIDTH_9_53_1": value  <=  8;
            "WIDTH_9_53_2": value  <=  8;
            "WIDTH_9_54_0": value  <=  6;
            "WIDTH_9_54_1": value  <=  3;
            "WIDTH_9_55_0": value  <=  10;
            "WIDTH_9_55_1": value  <=  5;
            "WIDTH_9_56_0": value  <=  2;
            "WIDTH_9_56_1": value  <=  1;
            "WIDTH_9_57_0": value  <=  6;
            "WIDTH_9_57_1": value  <=  3;
            "WIDTH_9_57_2": value  <=  3;
            "WIDTH_9_58_0": value  <=  8;
            "WIDTH_9_58_1": value  <=  8;
            "WIDTH_9_59_0": value  <=  6;
            "WIDTH_9_59_1": value  <=  3;
            "WIDTH_9_59_2": value  <=  3;
            "WIDTH_9_60_0": value  <=  6;
            "WIDTH_9_60_1": value  <=  3;
            "WIDTH_9_60_2": value  <=  3;
            "WIDTH_9_61_0": value  <=  1;
            "WIDTH_9_61_1": value  <=  1;
            "WIDTH_9_62_0": value  <=  2;
            "WIDTH_9_62_1": value  <=  1;
            "WIDTH_9_63_0": value  <=  2;
            "WIDTH_9_63_1": value  <=  2;
            "WIDTH_9_64_0": value  <=  2;
            "WIDTH_9_64_1": value  <=  2;
            "WIDTH_9_65_0": value  <=  4;
            "WIDTH_9_65_1": value  <=  4;
            "WIDTH_9_66_0": value  <=  2;
            "WIDTH_9_66_1": value  <=  1;
            "WIDTH_9_66_2": value  <=  1;
            "WIDTH_9_67_0": value  <=  11;
            "WIDTH_9_67_1": value  <=  11;
            "WIDTH_9_68_0": value  <=  4;
            "WIDTH_9_68_1": value  <=  4;
            "WIDTH_9_69_0": value  <=  8;
            "WIDTH_9_69_1": value  <=  4;
            "WIDTH_9_70_0": value  <=  1;
            "WIDTH_9_70_1": value  <=  1;
            "WIDTH_10_0_0": value  <=  6;
            "WIDTH_10_0_1": value  <=  3;
            "WIDTH_10_1_0": value  <=  6;
            "WIDTH_10_1_1": value  <=  3;
            "WIDTH_10_1_2": value  <=  3;
            "WIDTH_10_2_0": value  <=  8;
            "WIDTH_10_2_1": value  <=  4;
            "WIDTH_10_2_2": value  <=  4;
            "WIDTH_10_3_0": value  <=  20;
            "WIDTH_10_3_1": value  <=  20;
            "WIDTH_10_4_0": value  <=  2;
            "WIDTH_10_4_1": value  <=  2;
            "WIDTH_10_5_0": value  <=  12;
            "WIDTH_10_5_1": value  <=  4;
            "WIDTH_10_6_0": value  <=  4;
            "WIDTH_10_6_1": value  <=  4;
            "WIDTH_10_7_0": value  <=  7;
            "WIDTH_10_7_1": value  <=  7;
            "WIDTH_10_8_0": value  <=  3;
            "WIDTH_10_8_1": value  <=  1;
            "WIDTH_10_9_0": value  <=  2;
            "WIDTH_10_9_1": value  <=  2;
            "WIDTH_10_10_0": value  <=  4;
            "WIDTH_10_10_1": value  <=  4;
            "WIDTH_10_11_0": value  <=  6;
            "WIDTH_10_11_1": value  <=  6;
            "WIDTH_10_12_0": value  <=  6;
            "WIDTH_10_12_1": value  <=  2;
            "WIDTH_10_13_0": value  <=  4;
            "WIDTH_10_13_1": value  <=  4;
            "WIDTH_10_14_0": value  <=  5;
            "WIDTH_10_14_1": value  <=  5;
            "WIDTH_10_15_0": value  <=  2;
            "WIDTH_10_15_1": value  <=  2;
            "WIDTH_10_16_0": value  <=  4;
            "WIDTH_10_16_1": value  <=  4;
            "WIDTH_10_17_0": value  <=  6;
            "WIDTH_10_17_1": value  <=  3;
            "WIDTH_10_17_2": value  <=  3;
            "WIDTH_10_18_0": value  <=  3;
            "WIDTH_10_18_1": value  <=  1;
            "WIDTH_10_19_0": value  <=  4;
            "WIDTH_10_19_1": value  <=  4;
            "WIDTH_10_20_0": value  <=  4;
            "WIDTH_10_20_1": value  <=  4;
            "WIDTH_10_21_0": value  <=  12;
            "WIDTH_10_21_1": value  <=  4;
            "WIDTH_10_22_0": value  <=  6;
            "WIDTH_10_22_1": value  <=  2;
            "WIDTH_10_23_0": value  <=  3;
            "WIDTH_10_23_1": value  <=  1;
            "WIDTH_10_24_0": value  <=  2;
            "WIDTH_10_24_1": value  <=  2;
            "WIDTH_10_25_0": value  <=  7;
            "WIDTH_10_25_1": value  <=  7;
            "WIDTH_10_26_0": value  <=  15;
            "WIDTH_10_26_1": value  <=  15;
            "WIDTH_10_27_0": value  <=  6;
            "WIDTH_10_27_1": value  <=  3;
            "WIDTH_10_28_0": value  <=  3;
            "WIDTH_10_28_1": value  <=  1;
            "WIDTH_10_29_0": value  <=  6;
            "WIDTH_10_29_1": value  <=  3;
            "WIDTH_10_30_0": value  <=  20;
            "WIDTH_10_30_1": value  <=  20;
            "WIDTH_10_31_0": value  <=  6;
            "WIDTH_10_31_1": value  <=  3;
            "WIDTH_10_32_0": value  <=  6;
            "WIDTH_10_32_1": value  <=  3;
            "WIDTH_10_33_0": value  <=  1;
            "WIDTH_10_33_1": value  <=  1;
            "WIDTH_10_34_0": value  <=  4;
            "WIDTH_10_34_1": value  <=  2;
            "WIDTH_10_35_0": value  <=  18;
            "WIDTH_10_35_1": value  <=  9;
            "WIDTH_10_35_2": value  <=  9;
            "WIDTH_10_36_0": value  <=  1;
            "WIDTH_10_36_1": value  <=  1;
            "WIDTH_10_37_0": value  <=  10;
            "WIDTH_10_37_1": value  <=  5;
            "WIDTH_10_37_2": value  <=  5;
            "WIDTH_10_38_0": value  <=  2;
            "WIDTH_10_38_1": value  <=  1;
            "WIDTH_10_39_0": value  <=  3;
            "WIDTH_10_39_1": value  <=  1;
            "WIDTH_10_40_0": value  <=  12;
            "WIDTH_10_40_1": value  <=  4;
            "WIDTH_10_41_0": value  <=  4;
            "WIDTH_10_41_1": value  <=  4;
            "WIDTH_10_42_0": value  <=  3;
            "WIDTH_10_42_1": value  <=  1;
            "WIDTH_10_43_0": value  <=  4;
            "WIDTH_10_43_1": value  <=  4;
            "WIDTH_10_44_0": value  <=  4;
            "WIDTH_10_44_1": value  <=  4;
            "WIDTH_10_45_0": value  <=  1;
            "WIDTH_10_45_1": value  <=  1;
            "WIDTH_10_46_0": value  <=  8;
            "WIDTH_10_46_1": value  <=  8;
            "WIDTH_10_47_0": value  <=  6;
            "WIDTH_10_47_1": value  <=  2;
            "WIDTH_10_48_0": value  <=  4;
            "WIDTH_10_48_1": value  <=  4;
            "WIDTH_10_49_0": value  <=  14;
            "WIDTH_10_49_1": value  <=  14;
            "WIDTH_10_50_0": value  <=  6;
            "WIDTH_10_50_1": value  <=  6;
            "WIDTH_10_51_0": value  <=  10;
            "WIDTH_10_51_1": value  <=  10;
            "WIDTH_10_52_0": value  <=  3;
            "WIDTH_10_52_1": value  <=  1;
            "WIDTH_10_53_0": value  <=  2;
            "WIDTH_10_53_1": value  <=  1;
            "WIDTH_10_54_0": value  <=  6;
            "WIDTH_10_54_1": value  <=  2;
            "WIDTH_10_55_0": value  <=  3;
            "WIDTH_10_55_1": value  <=  1;
            "WIDTH_10_56_0": value  <=  2;
            "WIDTH_10_56_1": value  <=  2;
            "WIDTH_10_57_0": value  <=  3;
            "WIDTH_10_57_1": value  <=  3;
            "WIDTH_10_58_0": value  <=  4;
            "WIDTH_10_58_1": value  <=  2;
            "WIDTH_10_58_2": value  <=  2;
            "WIDTH_10_59_0": value  <=  2;
            "WIDTH_10_59_1": value  <=  2;
            "WIDTH_10_60_0": value  <=  2;
            "WIDTH_10_60_1": value  <=  2;
            "WIDTH_10_61_0": value  <=  4;
            "WIDTH_10_61_1": value  <=  4;
            "WIDTH_10_62_0": value  <=  20;
            "WIDTH_10_62_1": value  <=  10;
            "WIDTH_10_63_0": value  <=  8;
            "WIDTH_10_63_1": value  <=  4;
            "WIDTH_10_64_0": value  <=  8;
            "WIDTH_10_64_1": value  <=  4;
            "WIDTH_10_65_0": value  <=  3;
            "WIDTH_10_65_1": value  <=  1;
            "WIDTH_10_66_0": value  <=  3;
            "WIDTH_10_66_1": value  <=  1;
            "WIDTH_10_67_0": value  <=  3;
            "WIDTH_10_67_1": value  <=  1;
            "WIDTH_10_68_0": value  <=  3;
            "WIDTH_10_68_1": value  <=  1;
            "WIDTH_10_69_0": value  <=  6;
            "WIDTH_10_69_1": value  <=  3;
            "WIDTH_10_70_0": value  <=  2;
            "WIDTH_10_70_1": value  <=  2;
            "WIDTH_10_71_0": value  <=  1;
            "WIDTH_10_71_1": value  <=  1;
            "WIDTH_10_72_0": value  <=  2;
            "WIDTH_10_72_1": value  <=  1;
            "WIDTH_10_72_2": value  <=  1;
            "WIDTH_10_73_0": value  <=  18;
            "WIDTH_10_73_1": value  <=  9;
            "WIDTH_10_73_2": value  <=  9;
            "WIDTH_10_74_0": value  <=  2;
            "WIDTH_10_74_1": value  <=  1;
            "WIDTH_10_74_2": value  <=  1;
            "WIDTH_10_75_0": value  <=  20;
            "WIDTH_10_75_1": value  <=  20;
            "WIDTH_10_76_0": value  <=  2;
            "WIDTH_10_76_1": value  <=  2;
            "WIDTH_10_77_0": value  <=  4;
            "WIDTH_10_77_1": value  <=  4;
            "WIDTH_10_78_0": value  <=  2;
            "WIDTH_10_78_1": value  <=  2;
            "WIDTH_10_79_0": value  <=  2;
            "WIDTH_10_79_1": value  <=  2;
            "WIDTH_11_0_0": value  <=  10;
            "WIDTH_11_0_1": value  <=  10;
            "WIDTH_11_1_0": value  <=  6;
            "WIDTH_11_1_1": value  <=  3;
            "WIDTH_11_1_2": value  <=  3;
            "WIDTH_11_2_0": value  <=  3;
            "WIDTH_11_2_1": value  <=  3;
            "WIDTH_11_3_0": value  <=  4;
            "WIDTH_11_3_1": value  <=  2;
            "WIDTH_11_3_2": value  <=  2;
            "WIDTH_11_4_0": value  <=  4;
            "WIDTH_11_4_1": value  <=  4;
            "WIDTH_11_5_0": value  <=  4;
            "WIDTH_11_5_1": value  <=  2;
            "WIDTH_11_6_0": value  <=  4;
            "WIDTH_11_6_1": value  <=  2;
            "WIDTH_11_6_2": value  <=  2;
            "WIDTH_11_7_0": value  <=  4;
            "WIDTH_11_7_1": value  <=  2;
            "WIDTH_11_8_0": value  <=  8;
            "WIDTH_11_8_1": value  <=  4;
            "WIDTH_11_9_0": value  <=  2;
            "WIDTH_11_9_1": value  <=  2;
            "WIDTH_11_10_0": value  <=  5;
            "WIDTH_11_10_1": value  <=  5;
            "WIDTH_11_11_0": value  <=  4;
            "WIDTH_11_11_1": value  <=  2;
            "WIDTH_11_12_0": value  <=  8;
            "WIDTH_11_12_1": value  <=  8;
            "WIDTH_11_13_0": value  <=  6;
            "WIDTH_11_13_1": value  <=  3;
            "WIDTH_11_14_0": value  <=  6;
            "WIDTH_11_14_1": value  <=  3;
            "WIDTH_11_15_0": value  <=  8;
            "WIDTH_11_15_1": value  <=  4;
            "WIDTH_11_16_0": value  <=  3;
            "WIDTH_11_16_1": value  <=  1;
            "WIDTH_11_17_0": value  <=  6;
            "WIDTH_11_17_1": value  <=  3;
            "WIDTH_11_18_0": value  <=  2;
            "WIDTH_11_18_1": value  <=  2;
            "WIDTH_11_19_0": value  <=  4;
            "WIDTH_11_19_1": value  <=  4;
            "WIDTH_11_20_0": value  <=  2;
            "WIDTH_11_20_1": value  <=  1;
            "WIDTH_11_21_0": value  <=  2;
            "WIDTH_11_21_1": value  <=  2;
            "WIDTH_11_22_0": value  <=  2;
            "WIDTH_11_22_1": value  <=  2;
            "WIDTH_11_23_0": value  <=  2;
            "WIDTH_11_23_1": value  <=  2;
            "WIDTH_11_24_0": value  <=  4;
            "WIDTH_11_24_1": value  <=  4;
            "WIDTH_11_25_0": value  <=  2;
            "WIDTH_11_25_1": value  <=  2;
            "WIDTH_11_26_0": value  <=  2;
            "WIDTH_11_26_1": value  <=  2;
            "WIDTH_11_27_0": value  <=  6;
            "WIDTH_11_27_1": value  <=  6;
            "WIDTH_11_28_0": value  <=  2;
            "WIDTH_11_28_1": value  <=  1;
            "WIDTH_11_29_0": value  <=  4;
            "WIDTH_11_29_1": value  <=  4;
            "WIDTH_11_30_0": value  <=  2;
            "WIDTH_11_30_1": value  <=  1;
            "WIDTH_11_31_0": value  <=  14;
            "WIDTH_11_31_1": value  <=  7;
            "WIDTH_11_31_2": value  <=  7;
            "WIDTH_11_32_0": value  <=  6;
            "WIDTH_11_32_1": value  <=  3;
            "WIDTH_11_32_2": value  <=  3;
            "WIDTH_11_33_0": value  <=  6;
            "WIDTH_11_33_1": value  <=  6;
            "WIDTH_11_34_0": value  <=  12;
            "WIDTH_11_34_1": value  <=  12;
            "WIDTH_11_35_0": value  <=  7;
            "WIDTH_11_35_1": value  <=  7;
            "WIDTH_11_36_0": value  <=  18;
            "WIDTH_11_36_1": value  <=  18;
            "WIDTH_11_37_0": value  <=  2;
            "WIDTH_11_37_1": value  <=  1;
            "WIDTH_11_38_0": value  <=  3;
            "WIDTH_11_38_1": value  <=  1;
            "WIDTH_11_39_0": value  <=  3;
            "WIDTH_11_39_1": value  <=  1;
            "WIDTH_11_40_0": value  <=  3;
            "WIDTH_11_40_1": value  <=  3;
            "WIDTH_11_41_0": value  <=  6;
            "WIDTH_11_41_1": value  <=  2;
            "WIDTH_11_42_0": value  <=  6;
            "WIDTH_11_42_1": value  <=  2;
            "WIDTH_11_43_0": value  <=  5;
            "WIDTH_11_43_1": value  <=  5;
            "WIDTH_11_44_0": value  <=  6;
            "WIDTH_11_44_1": value  <=  2;
            "WIDTH_11_45_0": value  <=  6;
            "WIDTH_11_45_1": value  <=  3;
            "WIDTH_11_46_0": value  <=  14;
            "WIDTH_11_46_1": value  <=  7;
            "WIDTH_11_46_2": value  <=  7;
            "WIDTH_11_47_0": value  <=  4;
            "WIDTH_11_47_1": value  <=  2;
            "WIDTH_11_48_0": value  <=  12;
            "WIDTH_11_48_1": value  <=  6;
            "WIDTH_11_48_2": value  <=  6;
            "WIDTH_11_49_0": value  <=  5;
            "WIDTH_11_49_1": value  <=  5;
            "WIDTH_11_50_0": value  <=  4;
            "WIDTH_11_50_1": value  <=  4;
            "WIDTH_11_51_0": value  <=  2;
            "WIDTH_11_51_1": value  <=  1;
            "WIDTH_11_52_0": value  <=  2;
            "WIDTH_11_52_1": value  <=  1;
            "WIDTH_11_53_0": value  <=  3;
            "WIDTH_11_53_1": value  <=  1;
            "WIDTH_11_54_0": value  <=  3;
            "WIDTH_11_54_1": value  <=  3;
            "WIDTH_11_55_0": value  <=  3;
            "WIDTH_11_55_1": value  <=  1;
            "WIDTH_11_56_0": value  <=  6;
            "WIDTH_11_56_1": value  <=  3;
            "WIDTH_11_56_2": value  <=  3;
            "WIDTH_11_57_0": value  <=  4;
            "WIDTH_11_57_1": value  <=  4;
            "WIDTH_11_58_0": value  <=  3;
            "WIDTH_11_58_1": value  <=  3;
            "WIDTH_11_59_0": value  <=  3;
            "WIDTH_11_59_1": value  <=  3;
            "WIDTH_11_60_0": value  <=  16;
            "WIDTH_11_60_1": value  <=  8;
            "WIDTH_11_60_2": value  <=  8;
            "WIDTH_11_61_0": value  <=  3;
            "WIDTH_11_61_1": value  <=  3;
            "WIDTH_11_62_0": value  <=  5;
            "WIDTH_11_62_1": value  <=  5;
            "WIDTH_11_63_0": value  <=  4;
            "WIDTH_11_63_1": value  <=  4;
            "WIDTH_11_64_0": value  <=  3;
            "WIDTH_11_64_1": value  <=  3;
            "WIDTH_11_65_0": value  <=  2;
            "WIDTH_11_65_1": value  <=  2;
            "WIDTH_11_66_0": value  <=  4;
            "WIDTH_11_66_1": value  <=  4;
            "WIDTH_11_67_0": value  <=  4;
            "WIDTH_11_67_1": value  <=  4;
            "WIDTH_11_68_0": value  <=  6;
            "WIDTH_11_68_1": value  <=  2;
            "WIDTH_11_69_0": value  <=  3;
            "WIDTH_11_69_1": value  <=  3;
            "WIDTH_11_70_0": value  <=  18;
            "WIDTH_11_70_1": value  <=  6;
            "WIDTH_11_71_0": value  <=  3;
            "WIDTH_11_71_1": value  <=  3;
            "WIDTH_11_72_0": value  <=  3;
            "WIDTH_11_72_1": value  <=  3;
            "WIDTH_11_73_0": value  <=  6;
            "WIDTH_11_73_1": value  <=  6;
            "WIDTH_11_74_0": value  <=  8;
            "WIDTH_11_74_1": value  <=  8;
            "WIDTH_11_75_0": value  <=  4;
            "WIDTH_11_75_1": value  <=  2;
            "WIDTH_11_76_0": value  <=  4;
            "WIDTH_11_76_1": value  <=  2;
            "WIDTH_11_77_0": value  <=  2;
            "WIDTH_11_77_1": value  <=  2;
            "WIDTH_11_78_0": value  <=  6;
            "WIDTH_11_78_1": value  <=  2;
            "WIDTH_11_79_0": value  <=  3;
            "WIDTH_11_79_1": value  <=  3;
            "WIDTH_11_80_0": value  <=  3;
            "WIDTH_11_80_1": value  <=  1;
            "WIDTH_11_81_0": value  <=  16;
            "WIDTH_11_81_1": value  <=  16;
            "WIDTH_11_82_0": value  <=  16;
            "WIDTH_11_82_1": value  <=  16;
            "WIDTH_11_83_0": value  <=  15;
            "WIDTH_11_83_1": value  <=  5;
            "WIDTH_11_84_0": value  <=  7;
            "WIDTH_11_84_1": value  <=  7;
            "WIDTH_11_85_0": value  <=  2;
            "WIDTH_11_85_1": value  <=  2;
            "WIDTH_11_86_0": value  <=  16;
            "WIDTH_11_86_1": value  <=  8;
            "WIDTH_11_86_2": value  <=  8;
            "WIDTH_11_87_0": value  <=  4;
            "WIDTH_11_87_1": value  <=  2;
            "WIDTH_11_87_2": value  <=  2;
            "WIDTH_11_88_0": value  <=  2;
            "WIDTH_11_88_1": value  <=  2;
            "WIDTH_11_89_0": value  <=  4;
            "WIDTH_11_89_1": value  <=  2;
            "WIDTH_11_89_2": value  <=  2;
            "WIDTH_11_90_0": value  <=  8;
            "WIDTH_11_90_1": value  <=  8;
            "WIDTH_11_91_0": value  <=  4;
            "WIDTH_11_91_1": value  <=  4;
            "WIDTH_11_92_0": value  <=  5;
            "WIDTH_11_92_1": value  <=  5;
            "WIDTH_11_93_0": value  <=  4;
            "WIDTH_11_93_1": value  <=  2;
            "WIDTH_11_94_0": value  <=  6;
            "WIDTH_11_94_1": value  <=  2;
            "WIDTH_11_95_0": value  <=  3;
            "WIDTH_11_95_1": value  <=  1;
            "WIDTH_11_96_0": value  <=  3;
            "WIDTH_11_96_1": value  <=  1;
            "WIDTH_11_97_0": value  <=  6;
            "WIDTH_11_97_1": value  <=  6;
            "WIDTH_11_98_0": value  <=  4;
            "WIDTH_11_98_1": value  <=  2;
            "WIDTH_11_99_0": value  <=  6;
            "WIDTH_11_99_1": value  <=  3;
            "WIDTH_11_100_0": value  <=  1;
            "WIDTH_11_100_1": value  <=  1;
            "WIDTH_11_101_0": value  <=  10;
            "WIDTH_11_101_1": value  <=  5;
            "WIDTH_11_101_2": value  <=  5;
            "WIDTH_11_102_0": value  <=  12;
            "WIDTH_11_102_1": value  <=  6;
            "WIDTH_11_102_2": value  <=  6;
            "WIDTH_12_0_0": value  <=  6;
            "WIDTH_12_0_1": value  <=  3;
            "WIDTH_12_1_0": value  <=  6;
            "WIDTH_12_1_1": value  <=  3;
            "WIDTH_12_1_2": value  <=  3;
            "WIDTH_12_2_0": value  <=  2;
            "WIDTH_12_2_1": value  <=  2;
            "WIDTH_12_3_0": value  <=  6;
            "WIDTH_12_3_1": value  <=  3;
            "WIDTH_12_3_2": value  <=  3;
            "WIDTH_12_4_0": value  <=  2;
            "WIDTH_12_4_1": value  <=  2;
            "WIDTH_12_5_0": value  <=  6;
            "WIDTH_12_5_1": value  <=  2;
            "WIDTH_12_6_0": value  <=  12;
            "WIDTH_12_6_1": value  <=  4;
            "WIDTH_12_7_0": value  <=  6;
            "WIDTH_12_7_1": value  <=  6;
            "WIDTH_12_8_0": value  <=  3;
            "WIDTH_12_8_1": value  <=  1;
            "WIDTH_12_9_0": value  <=  3;
            "WIDTH_12_9_1": value  <=  3;
            "WIDTH_12_10_0": value  <=  17;
            "WIDTH_12_10_1": value  <=  17;
            "WIDTH_12_11_0": value  <=  4;
            "WIDTH_12_11_1": value  <=  2;
            "WIDTH_12_12_0": value  <=  4;
            "WIDTH_12_12_1": value  <=  4;
            "WIDTH_12_13_0": value  <=  2;
            "WIDTH_12_13_1": value  <=  1;
            "WIDTH_12_14_0": value  <=  6;
            "WIDTH_12_14_1": value  <=  2;
            "WIDTH_12_15_0": value  <=  2;
            "WIDTH_12_15_1": value  <=  2;
            "WIDTH_12_16_0": value  <=  3;
            "WIDTH_12_16_1": value  <=  3;
            "WIDTH_12_17_0": value  <=  12;
            "WIDTH_12_17_1": value  <=  12;
            "WIDTH_12_18_0": value  <=  4;
            "WIDTH_12_18_1": value  <=  2;
            "WIDTH_12_19_0": value  <=  3;
            "WIDTH_12_19_1": value  <=  3;
            "WIDTH_12_20_0": value  <=  6;
            "WIDTH_12_20_1": value  <=  2;
            "WIDTH_12_21_0": value  <=  3;
            "WIDTH_12_21_1": value  <=  3;
            "WIDTH_12_22_0": value  <=  3;
            "WIDTH_12_22_1": value  <=  1;
            "WIDTH_12_23_0": value  <=  2;
            "WIDTH_12_23_1": value  <=  2;
            "WIDTH_12_24_0": value  <=  6;
            "WIDTH_12_24_1": value  <=  6;
            "WIDTH_12_25_0": value  <=  4;
            "WIDTH_12_25_1": value  <=  4;
            "WIDTH_12_26_0": value  <=  2;
            "WIDTH_12_26_1": value  <=  2;
            "WIDTH_12_27_0": value  <=  12;
            "WIDTH_12_27_1": value  <=  4;
            "WIDTH_12_28_0": value  <=  3;
            "WIDTH_12_28_1": value  <=  3;
            "WIDTH_12_29_0": value  <=  1;
            "WIDTH_12_29_1": value  <=  1;
            "WIDTH_12_30_0": value  <=  3;
            "WIDTH_12_30_1": value  <=  1;
            "WIDTH_12_31_0": value  <=  5;
            "WIDTH_12_31_1": value  <=  5;
            "WIDTH_12_32_0": value  <=  5;
            "WIDTH_12_32_1": value  <=  5;
            "WIDTH_12_33_0": value  <=  2;
            "WIDTH_12_33_1": value  <=  1;
            "WIDTH_12_33_2": value  <=  1;
            "WIDTH_12_34_0": value  <=  3;
            "WIDTH_12_34_1": value  <=  1;
            "WIDTH_12_35_0": value  <=  2;
            "WIDTH_12_35_1": value  <=  2;
            "WIDTH_12_36_0": value  <=  2;
            "WIDTH_12_36_1": value  <=  2;
            "WIDTH_12_37_0": value  <=  12;
            "WIDTH_12_37_1": value  <=  12;
            "WIDTH_12_38_0": value  <=  3;
            "WIDTH_12_38_1": value  <=  3;
            "WIDTH_12_39_0": value  <=  2;
            "WIDTH_12_39_1": value  <=  1;
            "WIDTH_12_39_2": value  <=  1;
            "WIDTH_12_40_0": value  <=  1;
            "WIDTH_12_40_1": value  <=  1;
            "WIDTH_12_41_0": value  <=  13;
            "WIDTH_12_41_1": value  <=  13;
            "WIDTH_12_42_0": value  <=  15;
            "WIDTH_12_42_1": value  <=  5;
            "WIDTH_12_43_0": value  <=  12;
            "WIDTH_12_43_1": value  <=  4;
            "WIDTH_12_44_0": value  <=  4;
            "WIDTH_12_44_1": value  <=  4;
            "WIDTH_12_45_0": value  <=  1;
            "WIDTH_12_45_1": value  <=  1;
            "WIDTH_12_46_0": value  <=  5;
            "WIDTH_12_46_1": value  <=  5;
            "WIDTH_12_47_0": value  <=  7;
            "WIDTH_12_47_1": value  <=  7;
            "WIDTH_12_48_0": value  <=  6;
            "WIDTH_12_48_1": value  <=  3;
            "WIDTH_12_48_2": value  <=  3;
            "WIDTH_12_49_0": value  <=  4;
            "WIDTH_12_49_1": value  <=  4;
            "WIDTH_12_50_0": value  <=  2;
            "WIDTH_12_50_1": value  <=  2;
            "WIDTH_12_51_0": value  <=  3;
            "WIDTH_12_51_1": value  <=  1;
            "WIDTH_12_52_0": value  <=  4;
            "WIDTH_12_52_1": value  <=  4;
            "WIDTH_12_53_0": value  <=  4;
            "WIDTH_12_53_1": value  <=  4;
            "WIDTH_12_54_0": value  <=  3;
            "WIDTH_12_54_1": value  <=  1;
            "WIDTH_12_55_0": value  <=  2;
            "WIDTH_12_55_1": value  <=  1;
            "WIDTH_12_55_2": value  <=  1;
            "WIDTH_12_56_0": value  <=  2;
            "WIDTH_12_56_1": value  <=  1;
            "WIDTH_12_56_2": value  <=  1;
            "WIDTH_12_57_0": value  <=  4;
            "WIDTH_12_57_1": value  <=  4;
            "WIDTH_12_58_0": value  <=  3;
            "WIDTH_12_58_1": value  <=  1;
            "WIDTH_12_59_0": value  <=  6;
            "WIDTH_12_59_1": value  <=  6;
            "WIDTH_12_60_0": value  <=  3;
            "WIDTH_12_60_1": value  <=  1;
            "WIDTH_12_61_0": value  <=  10;
            "WIDTH_12_61_1": value  <=  5;
            "WIDTH_12_61_2": value  <=  5;
            "WIDTH_12_62_0": value  <=  8;
            "WIDTH_12_62_1": value  <=  4;
            "WIDTH_12_62_2": value  <=  4;
            "WIDTH_12_63_0": value  <=  6;
            "WIDTH_12_63_1": value  <=  2;
            "WIDTH_12_64_0": value  <=  6;
            "WIDTH_12_64_1": value  <=  2;
            "WIDTH_12_65_0": value  <=  3;
            "WIDTH_12_65_1": value  <=  1;
            "WIDTH_12_66_0": value  <=  2;
            "WIDTH_12_66_1": value  <=  1;
            "WIDTH_12_67_0": value  <=  1;
            "WIDTH_12_67_1": value  <=  1;
            "WIDTH_12_68_0": value  <=  2;
            "WIDTH_12_68_1": value  <=  1;
            "WIDTH_12_68_2": value  <=  1;
            "WIDTH_12_69_0": value  <=  1;
            "WIDTH_12_69_1": value  <=  1;
            "WIDTH_12_70_0": value  <=  3;
            "WIDTH_12_70_1": value  <=  1;
            "WIDTH_12_71_0": value  <=  2;
            "WIDTH_12_71_1": value  <=  1;
            "WIDTH_12_72_0": value  <=  8;
            "WIDTH_12_72_1": value  <=  8;
            "WIDTH_12_73_0": value  <=  15;
            "WIDTH_12_73_1": value  <=  15;
            "WIDTH_12_74_0": value  <=  12;
            "WIDTH_12_74_1": value  <=  12;
            "WIDTH_12_75_0": value  <=  4;
            "WIDTH_12_75_1": value  <=  2;
            "WIDTH_12_76_0": value  <=  3;
            "WIDTH_12_76_1": value  <=  1;
            "WIDTH_12_77_0": value  <=  4;
            "WIDTH_12_77_1": value  <=  2;
            "WIDTH_12_78_0": value  <=  6;
            "WIDTH_12_78_1": value  <=  2;
            "WIDTH_12_79_0": value  <=  4;
            "WIDTH_12_79_1": value  <=  2;
            "WIDTH_12_80_0": value  <=  4;
            "WIDTH_12_80_1": value  <=  2;
            "WIDTH_12_81_0": value  <=  3;
            "WIDTH_12_81_1": value  <=  3;
            "WIDTH_12_82_0": value  <=  3;
            "WIDTH_12_82_1": value  <=  3;
            "WIDTH_12_83_0": value  <=  4;
            "WIDTH_12_83_1": value  <=  4;
            "WIDTH_12_84_0": value  <=  2;
            "WIDTH_12_84_1": value  <=  1;
            "WIDTH_12_84_2": value  <=  1;
            "WIDTH_12_85_0": value  <=  4;
            "WIDTH_12_85_1": value  <=  4;
            "WIDTH_12_86_0": value  <=  4;
            "WIDTH_12_86_1": value  <=  4;
            "WIDTH_12_87_0": value  <=  1;
            "WIDTH_12_87_1": value  <=  1;
            "WIDTH_12_88_0": value  <=  3;
            "WIDTH_12_88_1": value  <=  1;
            "WIDTH_12_89_0": value  <=  3;
            "WIDTH_12_89_1": value  <=  1;
            "WIDTH_12_90_0": value  <=  3;
            "WIDTH_12_90_1": value  <=  1;
            "WIDTH_12_91_0": value  <=  4;
            "WIDTH_12_91_1": value  <=  2;
            "WIDTH_12_92_0": value  <=  5;
            "WIDTH_12_92_1": value  <=  5;
            "WIDTH_12_93_0": value  <=  6;
            "WIDTH_12_93_1": value  <=  3;
            "WIDTH_12_94_0": value  <=  18;
            "WIDTH_12_94_1": value  <=  6;
            "WIDTH_12_95_0": value  <=  4;
            "WIDTH_12_95_1": value  <=  2;
            "WIDTH_12_96_0": value  <=  4;
            "WIDTH_12_96_1": value  <=  2;
            "WIDTH_12_97_0": value  <=  1;
            "WIDTH_12_97_1": value  <=  1;
            "WIDTH_12_98_0": value  <=  2;
            "WIDTH_12_98_1": value  <=  1;
            "WIDTH_12_99_0": value  <=  2;
            "WIDTH_12_99_1": value  <=  1;
            "WIDTH_12_99_2": value  <=  1;
            "WIDTH_12_100_0": value  <=  4;
            "WIDTH_12_100_1": value  <=  4;
            "WIDTH_12_101_0": value  <=  2;
            "WIDTH_12_101_1": value  <=  1;
            "WIDTH_12_101_2": value  <=  1;
            "WIDTH_12_102_0": value  <=  4;
            "WIDTH_12_102_1": value  <=  2;
            "WIDTH_12_102_2": value  <=  2;
            "WIDTH_12_103_0": value  <=  7;
            "WIDTH_12_103_1": value  <=  7;
            "WIDTH_12_104_0": value  <=  6;
            "WIDTH_12_104_1": value  <=  3;
            "WIDTH_12_104_2": value  <=  3;
            "WIDTH_12_105_0": value  <=  3;
            "WIDTH_12_105_1": value  <=  1;
            "WIDTH_12_106_0": value  <=  5;
            "WIDTH_12_106_1": value  <=  5;
            "WIDTH_12_107_0": value  <=  1;
            "WIDTH_12_107_1": value  <=  1;
            "WIDTH_12_108_0": value  <=  18;
            "WIDTH_12_108_1": value  <=  9;
            "WIDTH_12_108_2": value  <=  9;
            "WIDTH_12_109_0": value  <=  2;
            "WIDTH_12_109_1": value  <=  1;
            "WIDTH_12_110_0": value  <=  4;
            "WIDTH_12_110_1": value  <=  2;
            "WIDTH_13_0_0": value  <=  6;
            "WIDTH_13_0_1": value  <=  2;
            "WIDTH_13_1_0": value  <=  18;
            "WIDTH_13_1_1": value  <=  6;
            "WIDTH_13_2_0": value  <=  2;
            "WIDTH_13_2_1": value  <=  2;
            "WIDTH_13_3_0": value  <=  19;
            "WIDTH_13_3_1": value  <=  19;
            "WIDTH_13_4_0": value  <=  3;
            "WIDTH_13_4_1": value  <=  3;
            "WIDTH_13_5_0": value  <=  4;
            "WIDTH_13_5_1": value  <=  2;
            "WIDTH_13_5_2": value  <=  2;
            "WIDTH_13_6_0": value  <=  4;
            "WIDTH_13_6_1": value  <=  2;
            "WIDTH_13_6_2": value  <=  2;
            "WIDTH_13_7_0": value  <=  10;
            "WIDTH_13_7_1": value  <=  10;
            "WIDTH_13_8_0": value  <=  14;
            "WIDTH_13_8_1": value  <=  14;
            "WIDTH_13_9_0": value  <=  10;
            "WIDTH_13_9_1": value  <=  5;
            "WIDTH_13_9_2": value  <=  5;
            "WIDTH_13_10_0": value  <=  2;
            "WIDTH_13_10_1": value  <=  2;
            "WIDTH_13_11_0": value  <=  6;
            "WIDTH_13_11_1": value  <=  3;
            "WIDTH_13_12_0": value  <=  2;
            "WIDTH_13_12_1": value  <=  2;
            "WIDTH_13_13_0": value  <=  6;
            "WIDTH_13_13_1": value  <=  3;
            "WIDTH_13_14_0": value  <=  6;
            "WIDTH_13_14_1": value  <=  3;
            "WIDTH_13_15_0": value  <=  6;
            "WIDTH_13_15_1": value  <=  2;
            "WIDTH_13_16_0": value  <=  6;
            "WIDTH_13_16_1": value  <=  2;
            "WIDTH_13_17_0": value  <=  2;
            "WIDTH_13_17_1": value  <=  2;
            "WIDTH_13_18_0": value  <=  1;
            "WIDTH_13_18_1": value  <=  1;
            "WIDTH_13_19_0": value  <=  2;
            "WIDTH_13_19_1": value  <=  2;
            "WIDTH_13_20_0": value  <=  3;
            "WIDTH_13_20_1": value  <=  1;
            "WIDTH_13_21_0": value  <=  9;
            "WIDTH_13_21_1": value  <=  9;
            "WIDTH_13_22_0": value  <=  4;
            "WIDTH_13_22_1": value  <=  4;
            "WIDTH_13_23_0": value  <=  2;
            "WIDTH_13_23_1": value  <=  2;
            "WIDTH_13_24_0": value  <=  2;
            "WIDTH_13_24_1": value  <=  2;
            "WIDTH_13_25_0": value  <=  3;
            "WIDTH_13_25_1": value  <=  3;
            "WIDTH_13_26_0": value  <=  3;
            "WIDTH_13_26_1": value  <=  3;
            "WIDTH_13_27_0": value  <=  3;
            "WIDTH_13_27_1": value  <=  3;
            "WIDTH_13_28_0": value  <=  3;
            "WIDTH_13_28_1": value  <=  3;
            "WIDTH_13_29_0": value  <=  2;
            "WIDTH_13_29_1": value  <=  1;
            "WIDTH_13_30_0": value  <=  3;
            "WIDTH_13_30_1": value  <=  1;
            "WIDTH_13_31_0": value  <=  8;
            "WIDTH_13_31_1": value  <=  4;
            "WIDTH_13_31_2": value  <=  4;
            "WIDTH_13_32_0": value  <=  8;
            "WIDTH_13_32_1": value  <=  4;
            "WIDTH_13_32_2": value  <=  4;
            "WIDTH_13_33_0": value  <=  3;
            "WIDTH_13_33_1": value  <=  3;
            "WIDTH_13_34_0": value  <=  3;
            "WIDTH_13_34_1": value  <=  3;
            "WIDTH_13_35_0": value  <=  3;
            "WIDTH_13_35_1": value  <=  3;
            "WIDTH_13_36_0": value  <=  6;
            "WIDTH_13_36_1": value  <=  6;
            "WIDTH_13_37_0": value  <=  6;
            "WIDTH_13_37_1": value  <=  6;
            "WIDTH_13_38_0": value  <=  6;
            "WIDTH_13_38_1": value  <=  6;
            "WIDTH_13_39_0": value  <=  5;
            "WIDTH_13_39_1": value  <=  5;
            "WIDTH_13_40_0": value  <=  3;
            "WIDTH_13_40_1": value  <=  3;
            "WIDTH_13_41_0": value  <=  5;
            "WIDTH_13_41_1": value  <=  5;
            "WIDTH_13_42_0": value  <=  6;
            "WIDTH_13_42_1": value  <=  2;
            "WIDTH_13_43_0": value  <=  4;
            "WIDTH_13_43_1": value  <=  4;
            "WIDTH_13_44_0": value  <=  5;
            "WIDTH_13_44_1": value  <=  5;
            "WIDTH_13_45_0": value  <=  4;
            "WIDTH_13_45_1": value  <=  2;
            "WIDTH_13_45_2": value  <=  2;
            "WIDTH_13_46_0": value  <=  3;
            "WIDTH_13_46_1": value  <=  1;
            "WIDTH_13_47_0": value  <=  5;
            "WIDTH_13_47_1": value  <=  5;
            "WIDTH_13_48_0": value  <=  20;
            "WIDTH_13_48_1": value  <=  10;
            "WIDTH_13_48_2": value  <=  10;
            "WIDTH_13_49_0": value  <=  18;
            "WIDTH_13_49_1": value  <=  6;
            "WIDTH_13_50_0": value  <=  6;
            "WIDTH_13_50_1": value  <=  2;
            "WIDTH_13_51_0": value  <=  13;
            "WIDTH_13_51_1": value  <=  13;
            "WIDTH_13_52_0": value  <=  3;
            "WIDTH_13_52_1": value  <=  3;
            "WIDTH_13_53_0": value  <=  6;
            "WIDTH_13_53_1": value  <=  3;
            "WIDTH_13_53_2": value  <=  3;
            "WIDTH_13_54_0": value  <=  10;
            "WIDTH_13_54_1": value  <=  5;
            "WIDTH_13_54_2": value  <=  5;
            "WIDTH_13_55_0": value  <=  1;
            "WIDTH_13_55_1": value  <=  1;
            "WIDTH_13_56_0": value  <=  4;
            "WIDTH_13_56_1": value  <=  4;
            "WIDTH_13_57_0": value  <=  2;
            "WIDTH_13_57_1": value  <=  2;
            "WIDTH_13_58_0": value  <=  2;
            "WIDTH_13_58_1": value  <=  2;
            "WIDTH_13_59_0": value  <=  9;
            "WIDTH_13_59_1": value  <=  9;
            "WIDTH_13_60_0": value  <=  2;
            "WIDTH_13_60_1": value  <=  2;
            "WIDTH_13_61_0": value  <=  3;
            "WIDTH_13_61_1": value  <=  3;
            "WIDTH_13_62_0": value  <=  9;
            "WIDTH_13_62_1": value  <=  9;
            "WIDTH_13_63_0": value  <=  3;
            "WIDTH_13_63_1": value  <=  3;
            "WIDTH_13_64_0": value  <=  3;
            "WIDTH_13_64_1": value  <=  3;
            "WIDTH_13_65_0": value  <=  11;
            "WIDTH_13_65_1": value  <=  11;
            "WIDTH_13_66_0": value  <=  5;
            "WIDTH_13_66_1": value  <=  5;
            "WIDTH_13_67_0": value  <=  18;
            "WIDTH_13_67_1": value  <=  18;
            "WIDTH_13_68_0": value  <=  5;
            "WIDTH_13_68_1": value  <=  5;
            "WIDTH_13_69_0": value  <=  12;
            "WIDTH_13_69_1": value  <=  4;
            "WIDTH_13_70_0": value  <=  6;
            "WIDTH_13_70_1": value  <=  3;
            "WIDTH_13_70_2": value  <=  3;
            "WIDTH_13_71_0": value  <=  12;
            "WIDTH_13_71_1": value  <=  4;
            "WIDTH_13_72_0": value  <=  12;
            "WIDTH_13_72_1": value  <=  4;
            "WIDTH_13_73_0": value  <=  6;
            "WIDTH_13_73_1": value  <=  3;
            "WIDTH_13_74_0": value  <=  16;
            "WIDTH_13_74_1": value  <=  16;
            "WIDTH_13_75_0": value  <=  10;
            "WIDTH_13_75_1": value  <=  10;
            "WIDTH_13_76_0": value  <=  10;
            "WIDTH_13_76_1": value  <=  5;
            "WIDTH_13_77_0": value  <=  2;
            "WIDTH_13_77_1": value  <=  2;
            "WIDTH_13_78_0": value  <=  2;
            "WIDTH_13_78_1": value  <=  2;
            "WIDTH_13_79_0": value  <=  3;
            "WIDTH_13_79_1": value  <=  1;
            "WIDTH_13_80_0": value  <=  4;
            "WIDTH_13_80_1": value  <=  2;
            "WIDTH_13_81_0": value  <=  6;
            "WIDTH_13_81_1": value  <=  2;
            "WIDTH_13_82_0": value  <=  12;
            "WIDTH_13_82_1": value  <=  6;
            "WIDTH_13_82_2": value  <=  6;
            "WIDTH_13_83_0": value  <=  6;
            "WIDTH_13_83_1": value  <=  2;
            "WIDTH_13_84_0": value  <=  6;
            "WIDTH_13_84_1": value  <=  2;
            "WIDTH_13_85_0": value  <=  6;
            "WIDTH_13_85_1": value  <=  3;
            "WIDTH_13_86_0": value  <=  6;
            "WIDTH_13_86_1": value  <=  3;
            "WIDTH_13_87_0": value  <=  6;
            "WIDTH_13_87_1": value  <=  2;
            "WIDTH_13_88_0": value  <=  6;
            "WIDTH_13_88_1": value  <=  2;
            "WIDTH_13_89_0": value  <=  3;
            "WIDTH_13_89_1": value  <=  3;
            "WIDTH_13_90_0": value  <=  6;
            "WIDTH_13_90_1": value  <=  2;
            "WIDTH_13_91_0": value  <=  18;
            "WIDTH_13_91_1": value  <=  9;
            "WIDTH_13_91_2": value  <=  9;
            "WIDTH_13_92_0": value  <=  10;
            "WIDTH_13_92_1": value  <=  10;
            "WIDTH_13_93_0": value  <=  4;
            "WIDTH_13_93_1": value  <=  4;
            "WIDTH_13_94_0": value  <=  3;
            "WIDTH_13_94_1": value  <=  3;
            "WIDTH_13_95_0": value  <=  16;
            "WIDTH_13_95_1": value  <=  16;
            "WIDTH_13_96_0": value  <=  12;
            "WIDTH_13_96_1": value  <=  6;
            "WIDTH_13_96_2": value  <=  6;
            "WIDTH_13_97_0": value  <=  2;
            "WIDTH_13_97_1": value  <=  1;
            "WIDTH_13_97_2": value  <=  1;
            "WIDTH_13_98_0": value  <=  10;
            "WIDTH_13_98_1": value  <=  5;
            "WIDTH_13_98_2": value  <=  5;
            "WIDTH_13_99_0": value  <=  3;
            "WIDTH_13_99_1": value  <=  3;
            "WIDTH_13_100_0": value  <=  9;
            "WIDTH_13_100_1": value  <=  9;
            "WIDTH_13_101_0": value  <=  2;
            "WIDTH_13_101_1": value  <=  2;
            "WIDTH_14_0_0": value  <=  13;
            "WIDTH_14_0_1": value  <=  13;
            "WIDTH_14_1_0": value  <=  6;
            "WIDTH_14_1_1": value  <=  3;
            "WIDTH_14_1_2": value  <=  3;
            "WIDTH_14_2_0": value  <=  6;
            "WIDTH_14_2_1": value  <=  3;
            "WIDTH_14_3_0": value  <=  2;
            "WIDTH_14_3_1": value  <=  2;
            "WIDTH_14_4_0": value  <=  3;
            "WIDTH_14_4_1": value  <=  3;
            "WIDTH_14_5_0": value  <=  8;
            "WIDTH_14_5_1": value  <=  8;
            "WIDTH_14_6_0": value  <=  10;
            "WIDTH_14_6_1": value  <=  10;
            "WIDTH_14_7_0": value  <=  3;
            "WIDTH_14_7_1": value  <=  3;
            "WIDTH_14_8_0": value  <=  4;
            "WIDTH_14_8_1": value  <=  2;
            "WIDTH_14_9_0": value  <=  3;
            "WIDTH_14_9_1": value  <=  3;
            "WIDTH_14_10_0": value  <=  8;
            "WIDTH_14_10_1": value  <=  8;
            "WIDTH_14_11_0": value  <=  6;
            "WIDTH_14_11_1": value  <=  6;
            "WIDTH_14_12_0": value  <=  3;
            "WIDTH_14_12_1": value  <=  3;
            "WIDTH_14_13_0": value  <=  3;
            "WIDTH_14_13_1": value  <=  3;
            "WIDTH_14_14_0": value  <=  4;
            "WIDTH_14_14_1": value  <=  2;
            "WIDTH_14_14_2": value  <=  2;
            "WIDTH_14_15_0": value  <=  3;
            "WIDTH_14_15_1": value  <=  3;
            "WIDTH_14_16_0": value  <=  4;
            "WIDTH_14_16_1": value  <=  4;
            "WIDTH_14_17_0": value  <=  6;
            "WIDTH_14_17_1": value  <=  3;
            "WIDTH_14_17_2": value  <=  3;
            "WIDTH_14_18_0": value  <=  3;
            "WIDTH_14_18_1": value  <=  1;
            "WIDTH_14_19_0": value  <=  4;
            "WIDTH_14_19_1": value  <=  4;
            "WIDTH_14_20_0": value  <=  8;
            "WIDTH_14_20_1": value  <=  4;
            "WIDTH_14_20_2": value  <=  4;
            "WIDTH_14_21_0": value  <=  2;
            "WIDTH_14_21_1": value  <=  1;
            "WIDTH_14_21_2": value  <=  1;
            "WIDTH_14_22_0": value  <=  8;
            "WIDTH_14_22_1": value  <=  4;
            "WIDTH_14_22_2": value  <=  4;
            "WIDTH_14_23_0": value  <=  6;
            "WIDTH_14_23_1": value  <=  3;
            "WIDTH_14_23_2": value  <=  3;
            "WIDTH_14_24_0": value  <=  1;
            "WIDTH_14_24_1": value  <=  1;
            "WIDTH_14_25_0": value  <=  4;
            "WIDTH_14_25_1": value  <=  4;
            "WIDTH_14_26_0": value  <=  2;
            "WIDTH_14_26_1": value  <=  2;
            "WIDTH_14_27_0": value  <=  14;
            "WIDTH_14_27_1": value  <=  7;
            "WIDTH_14_27_2": value  <=  7;
            "WIDTH_14_28_0": value  <=  4;
            "WIDTH_14_28_1": value  <=  4;
            "WIDTH_14_29_0": value  <=  6;
            "WIDTH_14_29_1": value  <=  2;
            "WIDTH_14_30_0": value  <=  6;
            "WIDTH_14_30_1": value  <=  2;
            "WIDTH_14_31_0": value  <=  16;
            "WIDTH_14_31_1": value  <=  16;
            "WIDTH_14_32_0": value  <=  4;
            "WIDTH_14_32_1": value  <=  2;
            "WIDTH_14_33_0": value  <=  12;
            "WIDTH_14_33_1": value  <=  6;
            "WIDTH_14_33_2": value  <=  6;
            "WIDTH_14_34_0": value  <=  3;
            "WIDTH_14_34_1": value  <=  1;
            "WIDTH_14_35_0": value  <=  4;
            "WIDTH_14_35_1": value  <=  2;
            "WIDTH_14_35_2": value  <=  2;
            "WIDTH_14_36_0": value  <=  4;
            "WIDTH_14_36_1": value  <=  4;
            "WIDTH_14_37_0": value  <=  3;
            "WIDTH_14_37_1": value  <=  1;
            "WIDTH_14_38_0": value  <=  3;
            "WIDTH_14_38_1": value  <=  3;
            "WIDTH_14_39_0": value  <=  9;
            "WIDTH_14_39_1": value  <=  3;
            "WIDTH_14_40_0": value  <=  2;
            "WIDTH_14_40_1": value  <=  1;
            "WIDTH_14_41_0": value  <=  2;
            "WIDTH_14_41_1": value  <=  2;
            "WIDTH_14_42_0": value  <=  4;
            "WIDTH_14_42_1": value  <=  4;
            "WIDTH_14_43_0": value  <=  8;
            "WIDTH_14_43_1": value  <=  8;
            "WIDTH_14_44_0": value  <=  7;
            "WIDTH_14_44_1": value  <=  7;
            "WIDTH_14_45_0": value  <=  8;
            "WIDTH_14_45_1": value  <=  8;
            "WIDTH_14_46_0": value  <=  3;
            "WIDTH_14_46_1": value  <=  1;
            "WIDTH_14_47_0": value  <=  6;
            "WIDTH_14_47_1": value  <=  3;
            "WIDTH_14_47_2": value  <=  3;
            "WIDTH_14_48_0": value  <=  6;
            "WIDTH_14_48_1": value  <=  3;
            "WIDTH_14_48_2": value  <=  3;
            "WIDTH_14_49_0": value  <=  18;
            "WIDTH_14_49_1": value  <=  9;
            "WIDTH_14_49_2": value  <=  9;
            "WIDTH_14_50_0": value  <=  2;
            "WIDTH_14_50_1": value  <=  1;
            "WIDTH_14_51_0": value  <=  4;
            "WIDTH_14_51_1": value  <=  2;
            "WIDTH_14_51_2": value  <=  2;
            "WIDTH_14_52_0": value  <=  3;
            "WIDTH_14_52_1": value  <=  3;
            "WIDTH_14_53_0": value  <=  1;
            "WIDTH_14_53_1": value  <=  1;
            "WIDTH_14_54_0": value  <=  5;
            "WIDTH_14_54_1": value  <=  5;
            "WIDTH_14_55_0": value  <=  4;
            "WIDTH_14_55_1": value  <=  2;
            "WIDTH_14_55_2": value  <=  2;
            "WIDTH_14_56_0": value  <=  4;
            "WIDTH_14_56_1": value  <=  2;
            "WIDTH_14_56_2": value  <=  2;
            "WIDTH_14_57_0": value  <=  1;
            "WIDTH_14_57_1": value  <=  1;
            "WIDTH_14_58_0": value  <=  2;
            "WIDTH_14_58_1": value  <=  2;
            "WIDTH_14_59_0": value  <=  2;
            "WIDTH_14_59_1": value  <=  1;
            "WIDTH_14_60_0": value  <=  2;
            "WIDTH_14_60_1": value  <=  1;
            "WIDTH_14_61_0": value  <=  3;
            "WIDTH_14_61_1": value  <=  3;
            "WIDTH_14_62_0": value  <=  4;
            "WIDTH_14_62_1": value  <=  2;
            "WIDTH_14_62_2": value  <=  2;
            "WIDTH_14_63_0": value  <=  2;
            "WIDTH_14_63_1": value  <=  2;
            "WIDTH_14_64_0": value  <=  9;
            "WIDTH_14_64_1": value  <=  9;
            "WIDTH_14_65_0": value  <=  2;
            "WIDTH_14_65_1": value  <=  2;
            "WIDTH_14_66_0": value  <=  2;
            "WIDTH_14_66_1": value  <=  2;
            "WIDTH_14_67_0": value  <=  18;
            "WIDTH_14_67_1": value  <=  18;
            "WIDTH_14_68_0": value  <=  4;
            "WIDTH_14_68_1": value  <=  4;
            "WIDTH_14_69_0": value  <=  6;
            "WIDTH_14_69_1": value  <=  6;
            "WIDTH_14_70_0": value  <=  2;
            "WIDTH_14_70_1": value  <=  2;
            "WIDTH_14_71_0": value  <=  3;
            "WIDTH_14_71_1": value  <=  1;
            "WIDTH_14_72_0": value  <=  18;
            "WIDTH_14_72_1": value  <=  6;
            "WIDTH_14_73_0": value  <=  3;
            "WIDTH_14_73_1": value  <=  1;
            "WIDTH_14_74_0": value  <=  1;
            "WIDTH_14_74_1": value  <=  1;
            "WIDTH_14_75_0": value  <=  8;
            "WIDTH_14_75_1": value  <=  4;
            "WIDTH_14_76_0": value  <=  3;
            "WIDTH_14_76_1": value  <=  1;
            "WIDTH_14_77_0": value  <=  2;
            "WIDTH_14_77_1": value  <=  2;
            "WIDTH_14_78_0": value  <=  2;
            "WIDTH_14_78_1": value  <=  1;
            "WIDTH_14_78_2": value  <=  1;
            "WIDTH_14_79_0": value  <=  2;
            "WIDTH_14_79_1": value  <=  1;
            "WIDTH_14_80_0": value  <=  2;
            "WIDTH_14_80_1": value  <=  1;
            "WIDTH_14_81_0": value  <=  2;
            "WIDTH_14_81_1": value  <=  2;
            "WIDTH_14_82_0": value  <=  2;
            "WIDTH_14_82_1": value  <=  2;
            "WIDTH_14_83_0": value  <=  15;
            "WIDTH_14_83_1": value  <=  5;
            "WIDTH_14_84_0": value  <=  15;
            "WIDTH_14_84_1": value  <=  5;
            "WIDTH_14_85_0": value  <=  2;
            "WIDTH_14_85_1": value  <=  2;
            "WIDTH_14_86_0": value  <=  4;
            "WIDTH_14_86_1": value  <=  2;
            "WIDTH_14_87_0": value  <=  2;
            "WIDTH_14_87_1": value  <=  1;
            "WIDTH_14_88_0": value  <=  2;
            "WIDTH_14_88_1": value  <=  1;
            "WIDTH_14_89_0": value  <=  3;
            "WIDTH_14_89_1": value  <=  3;
            "WIDTH_14_90_0": value  <=  3;
            "WIDTH_14_90_1": value  <=  3;
            "WIDTH_14_91_0": value  <=  8;
            "WIDTH_14_91_1": value  <=  8;
            "WIDTH_14_92_0": value  <=  6;
            "WIDTH_14_92_1": value  <=  6;
            "WIDTH_14_93_0": value  <=  18;
            "WIDTH_14_93_1": value  <=  6;
            "WIDTH_14_94_0": value  <=  3;
            "WIDTH_14_94_1": value  <=  1;
            "WIDTH_14_95_0": value  <=  4;
            "WIDTH_14_95_1": value  <=  2;
            "WIDTH_14_95_2": value  <=  2;
            "WIDTH_14_96_0": value  <=  3;
            "WIDTH_14_96_1": value  <=  1;
            "WIDTH_14_97_0": value  <=  2;
            "WIDTH_14_97_1": value  <=  2;
            "WIDTH_14_98_0": value  <=  4;
            "WIDTH_14_98_1": value  <=  2;
            "WIDTH_14_98_2": value  <=  2;
            "WIDTH_14_99_0": value  <=  20;
            "WIDTH_14_99_1": value  <=  10;
            "WIDTH_14_99_2": value  <=  10;
            "WIDTH_14_100_0": value  <=  2;
            "WIDTH_14_100_1": value  <=  1;
            "WIDTH_14_101_0": value  <=  18;
            "WIDTH_14_101_1": value  <=  9;
            "WIDTH_14_101_2": value  <=  9;
            "WIDTH_14_102_0": value  <=  2;
            "WIDTH_14_102_1": value  <=  1;
            "WIDTH_14_103_0": value  <=  16;
            "WIDTH_14_103_1": value  <=  8;
            "WIDTH_14_103_2": value  <=  8;
            "WIDTH_14_104_0": value  <=  1;
            "WIDTH_14_104_1": value  <=  1;
            "WIDTH_14_105_0": value  <=  4;
            "WIDTH_14_105_1": value  <=  4;
            "WIDTH_14_106_0": value  <=  8;
            "WIDTH_14_106_1": value  <=  4;
            "WIDTH_14_106_2": value  <=  4;
            "WIDTH_14_107_0": value  <=  8;
            "WIDTH_14_107_1": value  <=  8;
            "WIDTH_14_108_0": value  <=  2;
            "WIDTH_14_108_1": value  <=  2;
            "WIDTH_14_109_0": value  <=  2;
            "WIDTH_14_109_1": value  <=  2;
            "WIDTH_14_110_0": value  <=  2;
            "WIDTH_14_110_1": value  <=  2;
            "WIDTH_14_111_0": value  <=  2;
            "WIDTH_14_111_1": value  <=  2;
            "WIDTH_14_112_0": value  <=  1;
            "WIDTH_14_112_1": value  <=  1;
            "WIDTH_14_113_0": value  <=  2;
            "WIDTH_14_113_1": value  <=  2;
            "WIDTH_14_114_0": value  <=  2;
            "WIDTH_14_114_1": value  <=  2;
            "WIDTH_14_115_0": value  <=  3;
            "WIDTH_14_115_1": value  <=  3;
            "WIDTH_14_116_0": value  <=  2;
            "WIDTH_14_116_1": value  <=  2;
            "WIDTH_14_117_0": value  <=  4;
            "WIDTH_14_117_1": value  <=  4;
            "WIDTH_14_118_0": value  <=  3;
            "WIDTH_14_118_1": value  <=  3;
            "WIDTH_14_119_0": value  <=  10;
            "WIDTH_14_119_1": value  <=  10;
            "WIDTH_14_120_0": value  <=  4;
            "WIDTH_14_120_1": value  <=  4;
            "WIDTH_14_121_0": value  <=  15;
            "WIDTH_14_121_1": value  <=  5;
            "WIDTH_14_122_0": value  <=  12;
            "WIDTH_14_122_1": value  <=  4;
            "WIDTH_14_123_0": value  <=  3;
            "WIDTH_14_123_1": value  <=  1;
            "WIDTH_14_124_0": value  <=  4;
            "WIDTH_14_124_1": value  <=  2;
            "WIDTH_14_125_0": value  <=  4;
            "WIDTH_14_125_1": value  <=  4;
            "WIDTH_14_126_0": value  <=  4;
            "WIDTH_14_126_1": value  <=  2;
            "WIDTH_14_127_0": value  <=  3;
            "WIDTH_14_127_1": value  <=  1;
            "WIDTH_14_128_0": value  <=  6;
            "WIDTH_14_128_1": value  <=  2;
            "WIDTH_14_129_0": value  <=  3;
            "WIDTH_14_129_1": value  <=  1;
            "WIDTH_14_130_0": value  <=  8;
            "WIDTH_14_130_1": value  <=  4;
            "WIDTH_14_131_0": value  <=  12;
            "WIDTH_14_131_1": value  <=  4;
            "WIDTH_14_132_0": value  <=  10;
            "WIDTH_14_132_1": value  <=  5;
            "WIDTH_14_133_0": value  <=  3;
            "WIDTH_14_133_1": value  <=  1;
            "WIDTH_14_134_0": value  <=  11;
            "WIDTH_14_134_1": value  <=  11;
            "WIDTH_15_0_0": value  <=  18;
            "WIDTH_15_0_1": value  <=  6;
            "WIDTH_15_1_0": value  <=  6;
            "WIDTH_15_1_1": value  <=  2;
            "WIDTH_15_2_0": value  <=  6;
            "WIDTH_15_2_1": value  <=  3;
            "WIDTH_15_2_2": value  <=  3;
            "WIDTH_15_3_0": value  <=  9;
            "WIDTH_15_3_1": value  <=  9;
            "WIDTH_15_4_0": value  <=  2;
            "WIDTH_15_4_1": value  <=  2;
            "WIDTH_15_5_0": value  <=  8;
            "WIDTH_15_5_1": value  <=  4;
            "WIDTH_15_5_2": value  <=  4;
            "WIDTH_15_6_0": value  <=  8;
            "WIDTH_15_6_1": value  <=  4;
            "WIDTH_15_6_2": value  <=  4;
            "WIDTH_15_7_0": value  <=  2;
            "WIDTH_15_7_1": value  <=  2;
            "WIDTH_15_8_0": value  <=  8;
            "WIDTH_15_8_1": value  <=  8;
            "WIDTH_15_9_0": value  <=  8;
            "WIDTH_15_9_1": value  <=  8;
            "WIDTH_15_10_0": value  <=  2;
            "WIDTH_15_10_1": value  <=  1;
            "WIDTH_15_10_2": value  <=  1;
            "WIDTH_15_11_0": value  <=  2;
            "WIDTH_15_11_1": value  <=  2;
            "WIDTH_15_12_0": value  <=  15;
            "WIDTH_15_12_1": value  <=  15;
            "WIDTH_15_13_0": value  <=  4;
            "WIDTH_15_13_1": value  <=  4;
            "WIDTH_15_14_0": value  <=  3;
            "WIDTH_15_14_1": value  <=  1;
            "WIDTH_15_15_0": value  <=  6;
            "WIDTH_15_15_1": value  <=  6;
            "WIDTH_15_16_0": value  <=  2;
            "WIDTH_15_16_1": value  <=  2;
            "WIDTH_15_17_0": value  <=  3;
            "WIDTH_15_17_1": value  <=  3;
            "WIDTH_15_18_0": value  <=  3;
            "WIDTH_15_18_1": value  <=  1;
            "WIDTH_15_19_0": value  <=  4;
            "WIDTH_15_19_1": value  <=  4;
            "WIDTH_15_20_0": value  <=  3;
            "WIDTH_15_20_1": value  <=  1;
            "WIDTH_15_21_0": value  <=  4;
            "WIDTH_15_21_1": value  <=  4;
            "WIDTH_15_22_0": value  <=  2;
            "WIDTH_15_22_1": value  <=  2;
            "WIDTH_15_23_0": value  <=  4;
            "WIDTH_15_23_1": value  <=  4;
            "WIDTH_15_24_0": value  <=  4;
            "WIDTH_15_24_1": value  <=  4;
            "WIDTH_15_25_0": value  <=  1;
            "WIDTH_15_25_1": value  <=  1;
            "WIDTH_15_26_0": value  <=  3;
            "WIDTH_15_26_1": value  <=  1;
            "WIDTH_15_27_0": value  <=  2;
            "WIDTH_15_27_1": value  <=  1;
            "WIDTH_15_27_2": value  <=  1;
            "WIDTH_15_28_0": value  <=  6;
            "WIDTH_15_28_1": value  <=  2;
            "WIDTH_15_29_0": value  <=  3;
            "WIDTH_15_29_1": value  <=  3;
            "WIDTH_15_30_0": value  <=  3;
            "WIDTH_15_30_1": value  <=  1;
            "WIDTH_15_31_0": value  <=  3;
            "WIDTH_15_31_1": value  <=  1;
            "WIDTH_15_32_0": value  <=  3;
            "WIDTH_15_32_1": value  <=  1;
            "WIDTH_15_33_0": value  <=  5;
            "WIDTH_15_33_1": value  <=  5;
            "WIDTH_15_34_0": value  <=  5;
            "WIDTH_15_34_1": value  <=  5;
            "WIDTH_15_35_0": value  <=  18;
            "WIDTH_15_35_1": value  <=  6;
            "WIDTH_15_36_0": value  <=  2;
            "WIDTH_15_36_1": value  <=  2;
            "WIDTH_15_37_0": value  <=  4;
            "WIDTH_15_37_1": value  <=  2;
            "WIDTH_15_37_2": value  <=  2;
            "WIDTH_15_38_0": value  <=  3;
            "WIDTH_15_38_1": value  <=  3;
            "WIDTH_15_39_0": value  <=  2;
            "WIDTH_15_39_1": value  <=  2;
            "WIDTH_15_40_0": value  <=  1;
            "WIDTH_15_40_1": value  <=  1;
            "WIDTH_15_41_0": value  <=  6;
            "WIDTH_15_41_1": value  <=  3;
            "WIDTH_15_42_0": value  <=  6;
            "WIDTH_15_42_1": value  <=  3;
            "WIDTH_15_43_0": value  <=  3;
            "WIDTH_15_43_1": value  <=  3;
            "WIDTH_15_44_0": value  <=  1;
            "WIDTH_15_44_1": value  <=  1;
            "WIDTH_15_45_0": value  <=  3;
            "WIDTH_15_45_1": value  <=  3;
            "WIDTH_15_46_0": value  <=  12;
            "WIDTH_15_46_1": value  <=  12;
            "WIDTH_15_47_0": value  <=  2;
            "WIDTH_15_47_1": value  <=  2;
            "WIDTH_15_48_0": value  <=  3;
            "WIDTH_15_48_1": value  <=  1;
            "WIDTH_15_49_0": value  <=  9;
            "WIDTH_15_49_1": value  <=  3;
            "WIDTH_15_50_0": value  <=  1;
            "WIDTH_15_50_1": value  <=  1;
            "WIDTH_15_51_0": value  <=  2;
            "WIDTH_15_51_1": value  <=  2;
            "WIDTH_15_52_0": value  <=  2;
            "WIDTH_15_52_1": value  <=  2;
            "WIDTH_15_53_0": value  <=  1;
            "WIDTH_15_53_1": value  <=  1;
            "WIDTH_15_54_0": value  <=  6;
            "WIDTH_15_54_1": value  <=  2;
            "WIDTH_15_55_0": value  <=  20;
            "WIDTH_15_55_1": value  <=  10;
            "WIDTH_15_56_0": value  <=  5;
            "WIDTH_15_56_1": value  <=  5;
            "WIDTH_15_57_0": value  <=  2;
            "WIDTH_15_57_1": value  <=  2;
            "WIDTH_15_58_0": value  <=  9;
            "WIDTH_15_58_1": value  <=  9;
            "WIDTH_15_59_0": value  <=  12;
            "WIDTH_15_59_1": value  <=  6;
            "WIDTH_15_59_2": value  <=  6;
            "WIDTH_15_60_0": value  <=  2;
            "WIDTH_15_60_1": value  <=  1;
            "WIDTH_15_61_0": value  <=  6;
            "WIDTH_15_61_1": value  <=  2;
            "WIDTH_15_62_0": value  <=  2;
            "WIDTH_15_62_1": value  <=  1;
            "WIDTH_15_62_2": value  <=  1;
            "WIDTH_15_63_0": value  <=  2;
            "WIDTH_15_63_1": value  <=  1;
            "WIDTH_15_64_0": value  <=  4;
            "WIDTH_15_64_1": value  <=  4;
            "WIDTH_15_65_0": value  <=  2;
            "WIDTH_15_65_1": value  <=  1;
            "WIDTH_15_66_0": value  <=  2;
            "WIDTH_15_66_1": value  <=  1;
            "WIDTH_15_67_0": value  <=  18;
            "WIDTH_15_67_1": value  <=  9;
            "WIDTH_15_67_2": value  <=  9;
            "WIDTH_15_68_0": value  <=  2;
            "WIDTH_15_68_1": value  <=  1;
            "WIDTH_15_68_2": value  <=  1;
            "WIDTH_15_69_0": value  <=  4;
            "WIDTH_15_69_1": value  <=  4;
            "WIDTH_15_70_0": value  <=  2;
            "WIDTH_15_70_1": value  <=  1;
            "WIDTH_15_70_2": value  <=  1;
            "WIDTH_15_71_0": value  <=  18;
            "WIDTH_15_71_1": value  <=  9;
            "WIDTH_15_71_2": value  <=  9;
            "WIDTH_15_72_0": value  <=  1;
            "WIDTH_15_72_1": value  <=  1;
            "WIDTH_15_73_0": value  <=  18;
            "WIDTH_15_73_1": value  <=  9;
            "WIDTH_15_73_2": value  <=  9;
            "WIDTH_15_74_0": value  <=  18;
            "WIDTH_15_74_1": value  <=  9;
            "WIDTH_15_74_2": value  <=  9;
            "WIDTH_15_75_0": value  <=  5;
            "WIDTH_15_75_1": value  <=  5;
            "WIDTH_15_76_0": value  <=  7;
            "WIDTH_15_76_1": value  <=  7;
            "WIDTH_15_77_0": value  <=  3;
            "WIDTH_15_77_1": value  <=  3;
            "WIDTH_15_78_0": value  <=  3;
            "WIDTH_15_78_1": value  <=  1;
            "WIDTH_15_79_0": value  <=  2;
            "WIDTH_15_79_1": value  <=  1;
            "WIDTH_15_80_0": value  <=  9;
            "WIDTH_15_80_1": value  <=  3;
            "WIDTH_15_81_0": value  <=  2;
            "WIDTH_15_81_1": value  <=  1;
            "WIDTH_15_81_2": value  <=  1;
            "WIDTH_15_82_0": value  <=  6;
            "WIDTH_15_82_1": value  <=  3;
            "WIDTH_15_82_2": value  <=  3;
            "WIDTH_15_83_0": value  <=  4;
            "WIDTH_15_83_1": value  <=  4;
            "WIDTH_15_84_0": value  <=  8;
            "WIDTH_15_84_1": value  <=  8;
            "WIDTH_15_85_0": value  <=  6;
            "WIDTH_15_85_1": value  <=  3;
            "WIDTH_15_86_0": value  <=  10;
            "WIDTH_15_86_1": value  <=  10;
            "WIDTH_15_87_0": value  <=  5;
            "WIDTH_15_87_1": value  <=  5;
            "WIDTH_15_88_0": value  <=  4;
            "WIDTH_15_88_1": value  <=  2;
            "WIDTH_15_88_2": value  <=  2;
            "WIDTH_15_89_0": value  <=  6;
            "WIDTH_15_89_1": value  <=  2;
            "WIDTH_15_90_0": value  <=  3;
            "WIDTH_15_90_1": value  <=  1;
            "WIDTH_15_91_0": value  <=  2;
            "WIDTH_15_91_1": value  <=  2;
            "WIDTH_15_92_0": value  <=  3;
            "WIDTH_15_92_1": value  <=  1;
            "WIDTH_15_93_0": value  <=  13;
            "WIDTH_15_93_1": value  <=  13;
            "WIDTH_15_94_0": value  <=  6;
            "WIDTH_15_94_1": value  <=  2;
            "WIDTH_15_95_0": value  <=  3;
            "WIDTH_15_95_1": value  <=  3;
            "WIDTH_15_96_0": value  <=  6;
            "WIDTH_15_96_1": value  <=  2;
            "WIDTH_15_97_0": value  <=  18;
            "WIDTH_15_97_1": value  <=  9;
            "WIDTH_15_97_2": value  <=  9;
            "WIDTH_15_98_0": value  <=  4;
            "WIDTH_15_98_1": value  <=  4;
            "WIDTH_15_99_0": value  <=  4;
            "WIDTH_15_99_1": value  <=  4;
            "WIDTH_15_100_0": value  <=  3;
            "WIDTH_15_100_1": value  <=  1;
            "WIDTH_15_101_0": value  <=  4;
            "WIDTH_15_101_1": value  <=  4;
            "WIDTH_15_102_0": value  <=  3;
            "WIDTH_15_102_1": value  <=  1;
            "WIDTH_15_103_0": value  <=  4;
            "WIDTH_15_103_1": value  <=  4;
            "WIDTH_15_104_0": value  <=  1;
            "WIDTH_15_104_1": value  <=  1;
            "WIDTH_15_105_0": value  <=  1;
            "WIDTH_15_105_1": value  <=  1;
            "WIDTH_15_106_0": value  <=  4;
            "WIDTH_15_106_1": value  <=  4;
            "WIDTH_15_107_0": value  <=  2;
            "WIDTH_15_107_1": value  <=  1;
            "WIDTH_15_107_2": value  <=  1;
            "WIDTH_15_108_0": value  <=  2;
            "WIDTH_15_108_1": value  <=  1;
            "WIDTH_15_108_2": value  <=  1;
            "WIDTH_15_109_0": value  <=  14;
            "WIDTH_15_109_1": value  <=  7;
            "WIDTH_15_109_2": value  <=  7;
            "WIDTH_15_110_0": value  <=  19;
            "WIDTH_15_110_1": value  <=  19;
            "WIDTH_15_111_0": value  <=  3;
            "WIDTH_15_111_1": value  <=  3;
            "WIDTH_15_112_0": value  <=  1;
            "WIDTH_15_112_1": value  <=  1;
            "WIDTH_15_113_0": value  <=  3;
            "WIDTH_15_113_1": value  <=  3;
            "WIDTH_15_114_0": value  <=  3;
            "WIDTH_15_114_1": value  <=  3;
            "WIDTH_15_115_0": value  <=  4;
            "WIDTH_15_115_1": value  <=  4;
            "WIDTH_15_116_0": value  <=  4;
            "WIDTH_15_116_1": value  <=  2;
            "WIDTH_15_117_0": value  <=  2;
            "WIDTH_15_117_1": value  <=  2;
            "WIDTH_15_118_0": value  <=  20;
            "WIDTH_15_118_1": value  <=  20;
            "WIDTH_15_119_0": value  <=  17;
            "WIDTH_15_119_1": value  <=  17;
            "WIDTH_15_120_0": value  <=  6;
            "WIDTH_15_120_1": value  <=  3;
            "WIDTH_15_120_2": value  <=  3;
            "WIDTH_15_121_0": value  <=  6;
            "WIDTH_15_121_1": value  <=  3;
            "WIDTH_15_122_0": value  <=  6;
            "WIDTH_15_122_1": value  <=  3;
            "WIDTH_15_123_0": value  <=  7;
            "WIDTH_15_123_1": value  <=  7;
            "WIDTH_15_124_0": value  <=  7;
            "WIDTH_15_124_1": value  <=  7;
            "WIDTH_15_125_0": value  <=  14;
            "WIDTH_15_125_1": value  <=  7;
            "WIDTH_15_125_2": value  <=  7;
            "WIDTH_15_126_0": value  <=  2;
            "WIDTH_15_126_1": value  <=  1;
            "WIDTH_15_126_2": value  <=  1;
            "WIDTH_15_127_0": value  <=  2;
            "WIDTH_15_127_1": value  <=  1;
            "WIDTH_15_128_0": value  <=  3;
            "WIDTH_15_128_1": value  <=  1;
            "WIDTH_15_129_0": value  <=  1;
            "WIDTH_15_129_1": value  <=  1;
            "WIDTH_15_130_0": value  <=  1;
            "WIDTH_15_130_1": value  <=  1;
            "WIDTH_15_131_0": value  <=  1;
            "WIDTH_15_131_1": value  <=  1;
            "WIDTH_15_132_0": value  <=  2;
            "WIDTH_15_132_1": value  <=  2;
            "WIDTH_15_133_0": value  <=  4;
            "WIDTH_15_133_1": value  <=  2;
            "WIDTH_15_133_2": value  <=  2;
            "WIDTH_15_134_0": value  <=  1;
            "WIDTH_15_134_1": value  <=  1;
            "WIDTH_15_135_0": value  <=  4;
            "WIDTH_15_135_1": value  <=  2;
            "WIDTH_15_136_0": value  <=  2;
            "WIDTH_15_136_1": value  <=  1;
            "WIDTH_15_136_2": value  <=  1;
            "WIDTH_16_0_0": value  <=  10;
            "WIDTH_16_0_1": value  <=  10;
            "WIDTH_16_1_0": value  <=  4;
            "WIDTH_16_1_1": value  <=  2;
            "WIDTH_16_2_0": value  <=  4;
            "WIDTH_16_2_1": value  <=  4;
            "WIDTH_16_3_0": value  <=  1;
            "WIDTH_16_3_1": value  <=  1;
            "WIDTH_16_4_0": value  <=  14;
            "WIDTH_16_4_1": value  <=  7;
            "WIDTH_16_4_2": value  <=  7;
            "WIDTH_16_5_0": value  <=  6;
            "WIDTH_16_5_1": value  <=  3;
            "WIDTH_16_5_2": value  <=  3;
            "WIDTH_16_6_0": value  <=  6;
            "WIDTH_16_6_1": value  <=  3;
            "WIDTH_16_6_2": value  <=  3;
            "WIDTH_16_7_0": value  <=  15;
            "WIDTH_16_7_1": value  <=  5;
            "WIDTH_16_8_0": value  <=  6;
            "WIDTH_16_8_1": value  <=  6;
            "WIDTH_16_9_0": value  <=  14;
            "WIDTH_16_9_1": value  <=  7;
            "WIDTH_16_9_2": value  <=  7;
            "WIDTH_16_10_0": value  <=  15;
            "WIDTH_16_10_1": value  <=  5;
            "WIDTH_16_11_0": value  <=  8;
            "WIDTH_16_11_1": value  <=  8;
            "WIDTH_16_12_0": value  <=  3;
            "WIDTH_16_12_1": value  <=  1;
            "WIDTH_16_13_0": value  <=  2;
            "WIDTH_16_13_1": value  <=  2;
            "WIDTH_16_14_0": value  <=  6;
            "WIDTH_16_14_1": value  <=  3;
            "WIDTH_16_14_2": value  <=  3;
            "WIDTH_16_15_0": value  <=  18;
            "WIDTH_16_15_1": value  <=  6;
            "WIDTH_16_16_0": value  <=  6;
            "WIDTH_16_16_1": value  <=  3;
            "WIDTH_16_17_0": value  <=  6;
            "WIDTH_16_17_1": value  <=  6;
            "WIDTH_16_18_0": value  <=  6;
            "WIDTH_16_18_1": value  <=  6;
            "WIDTH_16_19_0": value  <=  3;
            "WIDTH_16_19_1": value  <=  3;
            "WIDTH_16_20_0": value  <=  3;
            "WIDTH_16_20_1": value  <=  3;
            "WIDTH_16_21_0": value  <=  2;
            "WIDTH_16_21_1": value  <=  2;
            "WIDTH_16_22_0": value  <=  6;
            "WIDTH_16_22_1": value  <=  6;
            "WIDTH_16_23_0": value  <=  3;
            "WIDTH_16_23_1": value  <=  3;
            "WIDTH_16_24_0": value  <=  2;
            "WIDTH_16_24_1": value  <=  2;
            "WIDTH_16_25_0": value  <=  6;
            "WIDTH_16_25_1": value  <=  2;
            "WIDTH_16_26_0": value  <=  3;
            "WIDTH_16_26_1": value  <=  3;
            "WIDTH_16_27_0": value  <=  4;
            "WIDTH_16_27_1": value  <=  4;
            "WIDTH_16_28_0": value  <=  3;
            "WIDTH_16_28_1": value  <=  3;
            "WIDTH_16_29_0": value  <=  3;
            "WIDTH_16_29_1": value  <=  1;
            "WIDTH_16_30_0": value  <=  5;
            "WIDTH_16_30_1": value  <=  5;
            "WIDTH_16_31_0": value  <=  2;
            "WIDTH_16_31_1": value  <=  2;
            "WIDTH_16_32_0": value  <=  14;
            "WIDTH_16_32_1": value  <=  7;
            "WIDTH_16_33_0": value  <=  18;
            "WIDTH_16_33_1": value  <=  18;
            "WIDTH_16_34_0": value  <=  2;
            "WIDTH_16_34_1": value  <=  2;
            "WIDTH_16_35_0": value  <=  4;
            "WIDTH_16_35_1": value  <=  2;
            "WIDTH_16_35_2": value  <=  2;
            "WIDTH_16_36_0": value  <=  4;
            "WIDTH_16_36_1": value  <=  2;
            "WIDTH_16_36_2": value  <=  2;
            "WIDTH_16_37_0": value  <=  3;
            "WIDTH_16_37_1": value  <=  1;
            "WIDTH_16_38_0": value  <=  2;
            "WIDTH_16_38_1": value  <=  1;
            "WIDTH_16_39_0": value  <=  15;
            "WIDTH_16_39_1": value  <=  15;
            "WIDTH_16_40_0": value  <=  3;
            "WIDTH_16_40_1": value  <=  1;
            "WIDTH_16_41_0": value  <=  18;
            "WIDTH_16_41_1": value  <=  9;
            "WIDTH_16_41_2": value  <=  9;
            "WIDTH_16_42_0": value  <=  2;
            "WIDTH_16_42_1": value  <=  1;
            "WIDTH_16_43_0": value  <=  2;
            "WIDTH_16_43_1": value  <=  1;
            "WIDTH_16_44_0": value  <=  6;
            "WIDTH_16_44_1": value  <=  2;
            "WIDTH_16_45_0": value  <=  2;
            "WIDTH_16_45_1": value  <=  1;
            "WIDTH_16_46_0": value  <=  2;
            "WIDTH_16_46_1": value  <=  1;
            "WIDTH_16_47_0": value  <=  14;
            "WIDTH_16_47_1": value  <=  14;
            "WIDTH_16_48_0": value  <=  6;
            "WIDTH_16_48_1": value  <=  6;
            "WIDTH_16_49_0": value  <=  3;
            "WIDTH_16_49_1": value  <=  1;
            "WIDTH_16_50_0": value  <=  4;
            "WIDTH_16_50_1": value  <=  4;
            "WIDTH_16_51_0": value  <=  6;
            "WIDTH_16_51_1": value  <=  6;
            "WIDTH_16_52_0": value  <=  2;
            "WIDTH_16_52_1": value  <=  2;
            "WIDTH_16_53_0": value  <=  6;
            "WIDTH_16_53_1": value  <=  2;
            "WIDTH_16_54_0": value  <=  4;
            "WIDTH_16_54_1": value  <=  4;
            "WIDTH_16_55_0": value  <=  7;
            "WIDTH_16_55_1": value  <=  7;
            "WIDTH_16_56_0": value  <=  8;
            "WIDTH_16_56_1": value  <=  4;
            "WIDTH_16_56_2": value  <=  4;
            "WIDTH_16_57_0": value  <=  3;
            "WIDTH_16_57_1": value  <=  3;
            "WIDTH_16_58_0": value  <=  2;
            "WIDTH_16_58_1": value  <=  2;
            "WIDTH_16_59_0": value  <=  1;
            "WIDTH_16_59_1": value  <=  1;
            "WIDTH_16_60_0": value  <=  14;
            "WIDTH_16_60_1": value  <=  14;
            "WIDTH_16_61_0": value  <=  1;
            "WIDTH_16_61_1": value  <=  1;
            "WIDTH_16_62_0": value  <=  3;
            "WIDTH_16_62_1": value  <=  1;
            "WIDTH_16_63_0": value  <=  2;
            "WIDTH_16_63_1": value  <=  1;
            "WIDTH_16_64_0": value  <=  6;
            "WIDTH_16_64_1": value  <=  6;
            "WIDTH_16_65_0": value  <=  8;
            "WIDTH_16_65_1": value  <=  8;
            "WIDTH_16_66_0": value  <=  1;
            "WIDTH_16_66_1": value  <=  1;
            "WIDTH_16_67_0": value  <=  6;
            "WIDTH_16_67_1": value  <=  6;
            "WIDTH_16_68_0": value  <=  2;
            "WIDTH_16_68_1": value  <=  1;
            "WIDTH_16_69_0": value  <=  18;
            "WIDTH_16_69_1": value  <=  9;
            "WIDTH_16_69_2": value  <=  9;
            "WIDTH_16_70_0": value  <=  2;
            "WIDTH_16_70_1": value  <=  2;
            "WIDTH_16_71_0": value  <=  5;
            "WIDTH_16_71_1": value  <=  5;
            "WIDTH_16_72_0": value  <=  2;
            "WIDTH_16_72_1": value  <=  2;
            "WIDTH_16_73_0": value  <=  3;
            "WIDTH_16_73_1": value  <=  1;
            "WIDTH_16_74_0": value  <=  6;
            "WIDTH_16_74_1": value  <=  2;
            "WIDTH_16_75_0": value  <=  5;
            "WIDTH_16_75_1": value  <=  5;
            "WIDTH_16_76_0": value  <=  5;
            "WIDTH_16_76_1": value  <=  5;
            "WIDTH_16_77_0": value  <=  1;
            "WIDTH_16_77_1": value  <=  1;
            "WIDTH_16_78_0": value  <=  9;
            "WIDTH_16_78_1": value  <=  3;
            "WIDTH_16_79_0": value  <=  3;
            "WIDTH_16_79_1": value  <=  1;
            "WIDTH_16_80_0": value  <=  4;
            "WIDTH_16_80_1": value  <=  2;
            "WIDTH_16_81_0": value  <=  1;
            "WIDTH_16_81_1": value  <=  1;
            "WIDTH_16_82_0": value  <=  1;
            "WIDTH_16_82_1": value  <=  1;
            "WIDTH_16_83_0": value  <=  1;
            "WIDTH_16_83_1": value  <=  1;
            "WIDTH_16_84_0": value  <=  3;
            "WIDTH_16_84_1": value  <=  1;
            "WIDTH_16_85_0": value  <=  2;
            "WIDTH_16_85_1": value  <=  2;
            "WIDTH_16_86_0": value  <=  1;
            "WIDTH_16_86_1": value  <=  1;
            "WIDTH_16_87_0": value  <=  8;
            "WIDTH_16_87_1": value  <=  4;
            "WIDTH_16_87_2": value  <=  4;
            "WIDTH_16_88_0": value  <=  8;
            "WIDTH_16_88_1": value  <=  4;
            "WIDTH_16_88_2": value  <=  4;
            "WIDTH_16_89_0": value  <=  18;
            "WIDTH_16_89_1": value  <=  18;
            "WIDTH_16_90_0": value  <=  2;
            "WIDTH_16_90_1": value  <=  2;
            "WIDTH_16_91_0": value  <=  14;
            "WIDTH_16_91_1": value  <=  14;
            "WIDTH_16_92_0": value  <=  4;
            "WIDTH_16_92_1": value  <=  2;
            "WIDTH_16_93_0": value  <=  4;
            "WIDTH_16_93_1": value  <=  2;
            "WIDTH_16_93_2": value  <=  2;
            "WIDTH_16_94_0": value  <=  2;
            "WIDTH_16_94_1": value  <=  1;
            "WIDTH_16_94_2": value  <=  1;
            "WIDTH_16_95_0": value  <=  2;
            "WIDTH_16_95_1": value  <=  2;
            "WIDTH_16_96_0": value  <=  3;
            "WIDTH_16_96_1": value  <=  3;
            "WIDTH_16_97_0": value  <=  6;
            "WIDTH_16_97_1": value  <=  6;
            "WIDTH_16_98_0": value  <=  11;
            "WIDTH_16_98_1": value  <=  11;
            "WIDTH_16_99_0": value  <=  6;
            "WIDTH_16_99_1": value  <=  2;
            "WIDTH_16_100_0": value  <=  4;
            "WIDTH_16_100_1": value  <=  4;
            "WIDTH_16_101_0": value  <=  2;
            "WIDTH_16_101_1": value  <=  2;
            "WIDTH_16_102_0": value  <=  3;
            "WIDTH_16_102_1": value  <=  3;
            "WIDTH_16_103_0": value  <=  3;
            "WIDTH_16_103_1": value  <=  1;
            "WIDTH_16_104_0": value  <=  3;
            "WIDTH_16_104_1": value  <=  1;
            "WIDTH_16_105_0": value  <=  3;
            "WIDTH_16_105_1": value  <=  1;
            "WIDTH_16_106_0": value  <=  3;
            "WIDTH_16_106_1": value  <=  1;
            "WIDTH_16_107_0": value  <=  16;
            "WIDTH_16_107_1": value  <=  8;
            "WIDTH_16_107_2": value  <=  8;
            "WIDTH_16_108_0": value  <=  4;
            "WIDTH_16_108_1": value  <=  2;
            "WIDTH_16_109_0": value  <=  2;
            "WIDTH_16_109_1": value  <=  1;
            "WIDTH_16_110_0": value  <=  6;
            "WIDTH_16_110_1": value  <=  3;
            "WIDTH_16_111_0": value  <=  12;
            "WIDTH_16_111_1": value  <=  4;
            "WIDTH_16_112_0": value  <=  8;
            "WIDTH_16_112_1": value  <=  4;
            "WIDTH_16_112_2": value  <=  4;
            "WIDTH_16_113_0": value  <=  2;
            "WIDTH_16_113_1": value  <=  1;
            "WIDTH_16_113_2": value  <=  1;
            "WIDTH_16_114_0": value  <=  20;
            "WIDTH_16_114_1": value  <=  20;
            "WIDTH_16_115_0": value  <=  2;
            "WIDTH_16_115_1": value  <=  1;
            "WIDTH_16_116_0": value  <=  9;
            "WIDTH_16_116_1": value  <=  3;
            "WIDTH_16_117_0": value  <=  16;
            "WIDTH_16_117_1": value  <=  8;
            "WIDTH_16_118_0": value  <=  3;
            "WIDTH_16_118_1": value  <=  3;
            "WIDTH_16_119_0": value  <=  6;
            "WIDTH_16_119_1": value  <=  6;
            "WIDTH_16_120_0": value  <=  1;
            "WIDTH_16_120_1": value  <=  1;
            "WIDTH_16_121_0": value  <=  4;
            "WIDTH_16_121_1": value  <=  4;
            "WIDTH_16_122_0": value  <=  2;
            "WIDTH_16_122_1": value  <=  2;
            "WIDTH_16_123_0": value  <=  10;
            "WIDTH_16_123_1": value  <=  5;
            "WIDTH_16_124_0": value  <=  12;
            "WIDTH_16_124_1": value  <=  6;
            "WIDTH_16_125_0": value  <=  20;
            "WIDTH_16_125_1": value  <=  10;
            "WIDTH_16_125_2": value  <=  10;
            "WIDTH_16_126_0": value  <=  2;
            "WIDTH_16_126_1": value  <=  1;
            "WIDTH_16_126_2": value  <=  1;
            "WIDTH_16_127_0": value  <=  2;
            "WIDTH_16_127_1": value  <=  1;
            "WIDTH_16_127_2": value  <=  1;
            "WIDTH_16_128_0": value  <=  2;
            "WIDTH_16_128_1": value  <=  1;
            "WIDTH_16_128_2": value  <=  1;
            "WIDTH_16_129_0": value  <=  1;
            "WIDTH_16_129_1": value  <=  1;
            "WIDTH_16_130_0": value  <=  16;
            "WIDTH_16_130_1": value  <=  8;
            "WIDTH_16_130_2": value  <=  8;
            "WIDTH_16_131_0": value  <=  3;
            "WIDTH_16_131_1": value  <=  1;
            "WIDTH_16_132_0": value  <=  2;
            "WIDTH_16_132_1": value  <=  2;
            "WIDTH_16_133_0": value  <=  15;
            "WIDTH_16_133_1": value  <=  5;
            "WIDTH_16_134_0": value  <=  15;
            "WIDTH_16_134_1": value  <=  5;
            "WIDTH_16_135_0": value  <=  2;
            "WIDTH_16_135_1": value  <=  1;
            "WIDTH_16_136_0": value  <=  2;
            "WIDTH_16_136_1": value  <=  1;
            "WIDTH_16_137_0": value  <=  2;
            "WIDTH_16_137_1": value  <=  1;
            "WIDTH_16_138_0": value  <=  2;
            "WIDTH_16_138_1": value  <=  1;
            "WIDTH_16_139_0": value  <=  14;
            "WIDTH_16_139_1": value  <=  7;
            "WIDTH_17_0_0": value  <=  18;
            "WIDTH_17_0_1": value  <=  6;
            "WIDTH_17_1_0": value  <=  6;
            "WIDTH_17_1_1": value  <=  3;
            "WIDTH_17_1_2": value  <=  3;
            "WIDTH_17_2_0": value  <=  2;
            "WIDTH_17_2_1": value  <=  2;
            "WIDTH_17_3_0": value  <=  6;
            "WIDTH_17_3_1": value  <=  6;
            "WIDTH_17_4_0": value  <=  6;
            "WIDTH_17_4_1": value  <=  3;
            "WIDTH_17_4_2": value  <=  3;
            "WIDTH_17_5_0": value  <=  6;
            "WIDTH_17_5_1": value  <=  3;
            "WIDTH_17_5_2": value  <=  3;
            "WIDTH_17_6_0": value  <=  18;
            "WIDTH_17_6_1": value  <=  6;
            "WIDTH_17_7_0": value  <=  9;
            "WIDTH_17_7_1": value  <=  9;
            "WIDTH_17_8_0": value  <=  4;
            "WIDTH_17_8_1": value  <=  2;
            "WIDTH_17_9_0": value  <=  3;
            "WIDTH_17_9_1": value  <=  3;
            "WIDTH_17_10_0": value  <=  5;
            "WIDTH_17_10_1": value  <=  5;
            "WIDTH_17_11_0": value  <=  6;
            "WIDTH_17_11_1": value  <=  3;
            "WIDTH_17_11_2": value  <=  3;
            "WIDTH_17_12_0": value  <=  10;
            "WIDTH_17_12_1": value  <=  10;
            "WIDTH_17_13_0": value  <=  1;
            "WIDTH_17_13_1": value  <=  1;
            "WIDTH_17_14_0": value  <=  3;
            "WIDTH_17_14_1": value  <=  3;
            "WIDTH_17_15_0": value  <=  4;
            "WIDTH_17_15_1": value  <=  4;
            "WIDTH_17_16_0": value  <=  1;
            "WIDTH_17_16_1": value  <=  1;
            "WIDTH_17_17_0": value  <=  2;
            "WIDTH_17_17_1": value  <=  2;
            "WIDTH_17_18_0": value  <=  3;
            "WIDTH_17_18_1": value  <=  1;
            "WIDTH_17_19_0": value  <=  11;
            "WIDTH_17_19_1": value  <=  11;
            "WIDTH_17_20_0": value  <=  20;
            "WIDTH_17_20_1": value  <=  20;
            "WIDTH_17_21_0": value  <=  1;
            "WIDTH_17_21_1": value  <=  1;
            "WIDTH_17_22_0": value  <=  2;
            "WIDTH_17_22_1": value  <=  1;
            "WIDTH_17_23_0": value  <=  12;
            "WIDTH_17_23_1": value  <=  4;
            "WIDTH_17_24_0": value  <=  12;
            "WIDTH_17_24_1": value  <=  4;
            "WIDTH_17_25_0": value  <=  3;
            "WIDTH_17_25_1": value  <=  1;
            "WIDTH_17_26_0": value  <=  6;
            "WIDTH_17_26_1": value  <=  3;
            "WIDTH_17_27_0": value  <=  3;
            "WIDTH_17_27_1": value  <=  3;
            "WIDTH_17_28_0": value  <=  6;
            "WIDTH_17_28_1": value  <=  2;
            "WIDTH_17_29_0": value  <=  3;
            "WIDTH_17_29_1": value  <=  3;
            "WIDTH_17_30_0": value  <=  2;
            "WIDTH_17_30_1": value  <=  1;
            "WIDTH_17_31_0": value  <=  9;
            "WIDTH_17_31_1": value  <=  3;
            "WIDTH_17_32_0": value  <=  4;
            "WIDTH_17_32_1": value  <=  4;
            "WIDTH_17_33_0": value  <=  4;
            "WIDTH_17_33_1": value  <=  2;
            "WIDTH_17_34_0": value  <=  6;
            "WIDTH_17_34_1": value  <=  6;
            "WIDTH_17_35_0": value  <=  3;
            "WIDTH_17_35_1": value  <=  3;
            "WIDTH_17_36_0": value  <=  3;
            "WIDTH_17_36_1": value  <=  1;
            "WIDTH_17_37_0": value  <=  4;
            "WIDTH_17_37_1": value  <=  2;
            "WIDTH_17_38_0": value  <=  3;
            "WIDTH_17_38_1": value  <=  1;
            "WIDTH_17_39_0": value  <=  9;
            "WIDTH_17_39_1": value  <=  3;
            "WIDTH_17_40_0": value  <=  8;
            "WIDTH_17_40_1": value  <=  4;
            "WIDTH_17_40_2": value  <=  4;
            "WIDTH_17_41_0": value  <=  6;
            "WIDTH_17_41_1": value  <=  2;
            "WIDTH_17_42_0": value  <=  3;
            "WIDTH_17_42_1": value  <=  1;
            "WIDTH_17_43_0": value  <=  6;
            "WIDTH_17_43_1": value  <=  2;
            "WIDTH_17_44_0": value  <=  6;
            "WIDTH_17_44_1": value  <=  6;
            "WIDTH_17_45_0": value  <=  6;
            "WIDTH_17_45_1": value  <=  3;
            "WIDTH_17_45_2": value  <=  3;
            "WIDTH_17_46_0": value  <=  3;
            "WIDTH_17_46_1": value  <=  1;
            "WIDTH_17_47_0": value  <=  2;
            "WIDTH_17_47_1": value  <=  1;
            "WIDTH_17_47_2": value  <=  1;
            "WIDTH_17_48_0": value  <=  18;
            "WIDTH_17_48_1": value  <=  6;
            "WIDTH_17_49_0": value  <=  2;
            "WIDTH_17_49_1": value  <=  1;
            "WIDTH_17_49_2": value  <=  1;
            "WIDTH_17_50_0": value  <=  12;
            "WIDTH_17_50_1": value  <=  4;
            "WIDTH_17_51_0": value  <=  5;
            "WIDTH_17_51_1": value  <=  5;
            "WIDTH_17_52_0": value  <=  2;
            "WIDTH_17_52_1": value  <=  2;
            "WIDTH_17_53_0": value  <=  2;
            "WIDTH_17_53_1": value  <=  1;
            "WIDTH_17_54_0": value  <=  1;
            "WIDTH_17_54_1": value  <=  1;
            "WIDTH_17_55_0": value  <=  2;
            "WIDTH_17_55_1": value  <=  2;
            "WIDTH_17_56_0": value  <=  2;
            "WIDTH_17_56_1": value  <=  2;
            "WIDTH_17_57_0": value  <=  2;
            "WIDTH_17_57_1": value  <=  2;
            "WIDTH_17_58_0": value  <=  2;
            "WIDTH_17_58_1": value  <=  2;
            "WIDTH_17_59_0": value  <=  1;
            "WIDTH_17_59_1": value  <=  1;
            "WIDTH_17_60_0": value  <=  2;
            "WIDTH_17_60_1": value  <=  2;
            "WIDTH_17_61_0": value  <=  2;
            "WIDTH_17_61_1": value  <=  1;
            "WIDTH_17_61_2": value  <=  1;
            "WIDTH_17_62_0": value  <=  2;
            "WIDTH_17_62_1": value  <=  2;
            "WIDTH_17_63_0": value  <=  14;
            "WIDTH_17_63_1": value  <=  14;
            "WIDTH_17_64_0": value  <=  4;
            "WIDTH_17_64_1": value  <=  4;
            "WIDTH_17_65_0": value  <=  1;
            "WIDTH_17_65_1": value  <=  1;
            "WIDTH_17_66_0": value  <=  1;
            "WIDTH_17_66_1": value  <=  1;
            "WIDTH_17_67_0": value  <=  6;
            "WIDTH_17_67_1": value  <=  2;
            "WIDTH_17_68_0": value  <=  2;
            "WIDTH_17_68_1": value  <=  1;
            "WIDTH_17_68_2": value  <=  1;
            "WIDTH_17_69_0": value  <=  6;
            "WIDTH_17_69_1": value  <=  3;
            "WIDTH_17_69_2": value  <=  3;
            "WIDTH_17_70_0": value  <=  6;
            "WIDTH_17_70_1": value  <=  3;
            "WIDTH_17_70_2": value  <=  3;
            "WIDTH_17_71_0": value  <=  3;
            "WIDTH_17_71_1": value  <=  3;
            "WIDTH_17_72_0": value  <=  3;
            "WIDTH_17_72_1": value  <=  3;
            "WIDTH_17_73_0": value  <=  6;
            "WIDTH_17_73_1": value  <=  2;
            "WIDTH_17_74_0": value  <=  6;
            "WIDTH_17_74_1": value  <=  2;
            "WIDTH_17_75_0": value  <=  7;
            "WIDTH_17_75_1": value  <=  7;
            "WIDTH_17_76_0": value  <=  2;
            "WIDTH_17_76_1": value  <=  1;
            "WIDTH_17_76_2": value  <=  1;
            "WIDTH_17_77_0": value  <=  8;
            "WIDTH_17_77_1": value  <=  4;
            "WIDTH_17_77_2": value  <=  4;
            "WIDTH_17_78_0": value  <=  2;
            "WIDTH_17_78_1": value  <=  1;
            "WIDTH_17_78_2": value  <=  1;
            "WIDTH_17_79_0": value  <=  16;
            "WIDTH_17_79_1": value  <=  8;
            "WIDTH_17_79_2": value  <=  8;
            "WIDTH_17_80_0": value  <=  3;
            "WIDTH_17_80_1": value  <=  3;
            "WIDTH_17_81_0": value  <=  3;
            "WIDTH_17_81_1": value  <=  3;
            "WIDTH_17_82_0": value  <=  3;
            "WIDTH_17_82_1": value  <=  3;
            "WIDTH_17_83_0": value  <=  3;
            "WIDTH_17_83_1": value  <=  1;
            "WIDTH_17_84_0": value  <=  4;
            "WIDTH_17_84_1": value  <=  4;
            "WIDTH_17_85_0": value  <=  1;
            "WIDTH_17_85_1": value  <=  1;
            "WIDTH_17_86_0": value  <=  4;
            "WIDTH_17_86_1": value  <=  2;
            "WIDTH_17_86_2": value  <=  2;
            "WIDTH_17_87_0": value  <=  4;
            "WIDTH_17_87_1": value  <=  4;
            "WIDTH_17_88_0": value  <=  1;
            "WIDTH_17_88_1": value  <=  1;
            "WIDTH_17_89_0": value  <=  2;
            "WIDTH_17_89_1": value  <=  2;
            "WIDTH_17_90_0": value  <=  4;
            "WIDTH_17_90_1": value  <=  4;
            "WIDTH_17_91_0": value  <=  3;
            "WIDTH_17_91_1": value  <=  1;
            "WIDTH_17_92_0": value  <=  3;
            "WIDTH_17_92_1": value  <=  1;
            "WIDTH_17_93_0": value  <=  6;
            "WIDTH_17_93_1": value  <=  2;
            "WIDTH_17_94_0": value  <=  2;
            "WIDTH_17_94_1": value  <=  1;
            "WIDTH_17_95_0": value  <=  8;
            "WIDTH_17_95_1": value  <=  4;
            "WIDTH_17_95_2": value  <=  4;
            "WIDTH_17_96_0": value  <=  8;
            "WIDTH_17_96_1": value  <=  4;
            "WIDTH_17_96_2": value  <=  4;
            "WIDTH_17_97_0": value  <=  2;
            "WIDTH_17_97_1": value  <=  1;
            "WIDTH_17_97_2": value  <=  1;
            "WIDTH_17_98_0": value  <=  6;
            "WIDTH_17_98_1": value  <=  3;
            "WIDTH_17_99_0": value  <=  6;
            "WIDTH_17_99_1": value  <=  2;
            "WIDTH_17_100_0": value  <=  2;
            "WIDTH_17_100_1": value  <=  1;
            "WIDTH_17_100_2": value  <=  1;
            "WIDTH_17_101_0": value  <=  1;
            "WIDTH_17_101_1": value  <=  1;
            "WIDTH_17_102_0": value  <=  1;
            "WIDTH_17_102_1": value  <=  1;
            "WIDTH_17_103_0": value  <=  2;
            "WIDTH_17_103_1": value  <=  1;
            "WIDTH_17_104_0": value  <=  2;
            "WIDTH_17_104_1": value  <=  2;
            "WIDTH_17_105_0": value  <=  7;
            "WIDTH_17_105_1": value  <=  7;
            "WIDTH_17_106_0": value  <=  12;
            "WIDTH_17_106_1": value  <=  12;
            "WIDTH_17_107_0": value  <=  3;
            "WIDTH_17_107_1": value  <=  1;
            "WIDTH_17_108_0": value  <=  2;
            "WIDTH_17_108_1": value  <=  2;
            "WIDTH_17_109_0": value  <=  4;
            "WIDTH_17_109_1": value  <=  4;
            "WIDTH_17_110_0": value  <=  2;
            "WIDTH_17_110_1": value  <=  1;
            "WIDTH_17_110_2": value  <=  1;
            "WIDTH_17_111_0": value  <=  14;
            "WIDTH_17_111_1": value  <=  7;
            "WIDTH_17_111_2": value  <=  7;
            "WIDTH_17_112_0": value  <=  18;
            "WIDTH_17_112_1": value  <=  6;
            "WIDTH_17_113_0": value  <=  2;
            "WIDTH_17_113_1": value  <=  1;
            "WIDTH_17_113_2": value  <=  1;
            "WIDTH_17_114_0": value  <=  2;
            "WIDTH_17_114_1": value  <=  1;
            "WIDTH_17_114_2": value  <=  1;
            "WIDTH_17_115_0": value  <=  8;
            "WIDTH_17_115_1": value  <=  8;
            "WIDTH_17_116_0": value  <=  6;
            "WIDTH_17_116_1": value  <=  6;
            "WIDTH_17_117_0": value  <=  4;
            "WIDTH_17_117_1": value  <=  2;
            "WIDTH_17_117_2": value  <=  2;
            "WIDTH_17_118_0": value  <=  3;
            "WIDTH_17_118_1": value  <=  3;
            "WIDTH_17_119_0": value  <=  6;
            "WIDTH_17_119_1": value  <=  2;
            "WIDTH_17_120_0": value  <=  4;
            "WIDTH_17_120_1": value  <=  2;
            "WIDTH_17_121_0": value  <=  12;
            "WIDTH_17_121_1": value  <=  4;
            "WIDTH_17_122_0": value  <=  3;
            "WIDTH_17_122_1": value  <=  3;
            "WIDTH_17_123_0": value  <=  12;
            "WIDTH_17_123_1": value  <=  4;
            "WIDTH_17_124_0": value  <=  3;
            "WIDTH_17_124_1": value  <=  3;
            "WIDTH_17_125_0": value  <=  4;
            "WIDTH_17_125_1": value  <=  2;
            "WIDTH_17_126_0": value  <=  4;
            "WIDTH_17_126_1": value  <=  2;
            "WIDTH_17_127_0": value  <=  2;
            "WIDTH_17_127_1": value  <=  1;
            "WIDTH_17_127_2": value  <=  1;
            "WIDTH_17_128_0": value  <=  3;
            "WIDTH_17_128_1": value  <=  3;
            "WIDTH_17_129_0": value  <=  2;
            "WIDTH_17_129_1": value  <=  1;
            "WIDTH_17_129_2": value  <=  1;
            "WIDTH_17_130_0": value  <=  4;
            "WIDTH_17_130_1": value  <=  4;
            "WIDTH_17_131_0": value  <=  2;
            "WIDTH_17_131_1": value  <=  1;
            "WIDTH_17_131_2": value  <=  1;
            "WIDTH_17_132_0": value  <=  5;
            "WIDTH_17_132_1": value  <=  5;
            "WIDTH_17_133_0": value  <=  2;
            "WIDTH_17_133_1": value  <=  1;
            "WIDTH_17_133_2": value  <=  1;
            "WIDTH_17_134_0": value  <=  2;
            "WIDTH_17_134_1": value  <=  1;
            "WIDTH_17_134_2": value  <=  1;
            "WIDTH_17_135_0": value  <=  3;
            "WIDTH_17_135_1": value  <=  3;
            "WIDTH_17_136_0": value  <=  3;
            "WIDTH_17_136_1": value  <=  3;
            "WIDTH_17_137_0": value  <=  2;
            "WIDTH_17_137_1": value  <=  2;
            "WIDTH_17_138_0": value  <=  3;
            "WIDTH_17_138_1": value  <=  3;
            "WIDTH_17_139_0": value  <=  3;
            "WIDTH_17_139_1": value  <=  3;
            "WIDTH_17_140_0": value  <=  5;
            "WIDTH_17_140_1": value  <=  5;
            "WIDTH_17_141_0": value  <=  3;
            "WIDTH_17_141_1": value  <=  3;
            "WIDTH_17_142_0": value  <=  2;
            "WIDTH_17_142_1": value  <=  1;
            "WIDTH_17_142_2": value  <=  1;
            "WIDTH_17_143_0": value  <=  2;
            "WIDTH_17_143_1": value  <=  1;
            "WIDTH_17_143_2": value  <=  1;
            "WIDTH_17_144_0": value  <=  6;
            "WIDTH_17_144_1": value  <=  3;
            "WIDTH_17_145_0": value  <=  2;
            "WIDTH_17_145_1": value  <=  2;
            "WIDTH_17_146_0": value  <=  2;
            "WIDTH_17_146_1": value  <=  2;
            "WIDTH_17_147_0": value  <=  8;
            "WIDTH_17_147_1": value  <=  4;
            "WIDTH_17_148_0": value  <=  8;
            "WIDTH_17_148_1": value  <=  4;
            "WIDTH_17_149_0": value  <=  3;
            "WIDTH_17_149_1": value  <=  1;
            "WIDTH_17_150_0": value  <=  4;
            "WIDTH_17_150_1": value  <=  2;
            "WIDTH_17_151_0": value  <=  3;
            "WIDTH_17_151_1": value  <=  1;
            "WIDTH_17_152_0": value  <=  3;
            "WIDTH_17_152_1": value  <=  1;
            "WIDTH_17_153_0": value  <=  3;
            "WIDTH_17_153_1": value  <=  3;
            "WIDTH_17_154_0": value  <=  7;
            "WIDTH_17_154_1": value  <=  7;
            "WIDTH_17_155_0": value  <=  2;
            "WIDTH_17_155_1": value  <=  1;
            "WIDTH_17_155_2": value  <=  1;
            "WIDTH_17_156_0": value  <=  2;
            "WIDTH_17_156_1": value  <=  1;
            "WIDTH_17_156_2": value  <=  1;
            "WIDTH_17_157_0": value  <=  4;
            "WIDTH_17_157_1": value  <=  2;
            "WIDTH_17_157_2": value  <=  2;
            "WIDTH_17_158_0": value  <=  2;
            "WIDTH_17_158_1": value  <=  1;
            "WIDTH_17_158_2": value  <=  1;
            "WIDTH_17_159_0": value  <=  3;
            "WIDTH_17_159_1": value  <=  3;
            "WIDTH_18_0_0": value  <=  19;
            "WIDTH_18_0_1": value  <=  19;
            "WIDTH_18_1_0": value  <=  10;
            "WIDTH_18_1_1": value  <=  5;
            "WIDTH_18_2_0": value  <=  2;
            "WIDTH_18_2_1": value  <=  2;
            "WIDTH_18_3_0": value  <=  4;
            "WIDTH_18_3_1": value  <=  2;
            "WIDTH_18_4_0": value  <=  6;
            "WIDTH_18_4_1": value  <=  3;
            "WIDTH_18_4_2": value  <=  3;
            "WIDTH_18_5_0": value  <=  6;
            "WIDTH_18_5_1": value  <=  2;
            "WIDTH_18_6_0": value  <=  6;
            "WIDTH_18_6_1": value  <=  2;
            "WIDTH_18_7_0": value  <=  8;
            "WIDTH_18_7_1": value  <=  8;
            "WIDTH_18_8_0": value  <=  2;
            "WIDTH_18_8_1": value  <=  1;
            "WIDTH_18_9_0": value  <=  9;
            "WIDTH_18_9_1": value  <=  3;
            "WIDTH_18_10_0": value  <=  9;
            "WIDTH_18_10_1": value  <=  3;
            "WIDTH_18_11_0": value  <=  18;
            "WIDTH_18_11_1": value  <=  6;
            "WIDTH_18_12_0": value  <=  5;
            "WIDTH_18_12_1": value  <=  5;
            "WIDTH_18_13_0": value  <=  6;
            "WIDTH_18_13_1": value  <=  2;
            "WIDTH_18_14_0": value  <=  3;
            "WIDTH_18_14_1": value  <=  3;
            "WIDTH_18_15_0": value  <=  4;
            "WIDTH_18_15_1": value  <=  4;
            "WIDTH_18_16_0": value  <=  3;
            "WIDTH_18_16_1": value  <=  3;
            "WIDTH_18_17_0": value  <=  2;
            "WIDTH_18_17_1": value  <=  1;
            "WIDTH_18_18_0": value  <=  2;
            "WIDTH_18_18_1": value  <=  1;
            "WIDTH_18_19_0": value  <=  2;
            "WIDTH_18_19_1": value  <=  1;
            "WIDTH_18_20_0": value  <=  8;
            "WIDTH_18_20_1": value  <=  8;
            "WIDTH_18_21_0": value  <=  3;
            "WIDTH_18_21_1": value  <=  1;
            "WIDTH_18_22_0": value  <=  2;
            "WIDTH_18_22_1": value  <=  1;
            "WIDTH_18_23_0": value  <=  6;
            "WIDTH_18_23_1": value  <=  2;
            "WIDTH_18_24_0": value  <=  3;
            "WIDTH_18_24_1": value  <=  1;
            "WIDTH_18_25_0": value  <=  7;
            "WIDTH_18_25_1": value  <=  7;
            "WIDTH_18_26_0": value  <=  3;
            "WIDTH_18_26_1": value  <=  1;
            "WIDTH_18_27_0": value  <=  8;
            "WIDTH_18_27_1": value  <=  8;
            "WIDTH_18_28_0": value  <=  8;
            "WIDTH_18_28_1": value  <=  8;
            "WIDTH_18_29_0": value  <=  2;
            "WIDTH_18_29_1": value  <=  2;
            "WIDTH_18_30_0": value  <=  2;
            "WIDTH_18_30_1": value  <=  2;
            "WIDTH_18_31_0": value  <=  4;
            "WIDTH_18_31_1": value  <=  4;
            "WIDTH_18_32_0": value  <=  4;
            "WIDTH_18_32_1": value  <=  4;
            "WIDTH_18_33_0": value  <=  1;
            "WIDTH_18_33_1": value  <=  1;
            "WIDTH_18_34_0": value  <=  4;
            "WIDTH_18_34_1": value  <=  4;
            "WIDTH_18_35_0": value  <=  4;
            "WIDTH_18_35_1": value  <=  2;
            "WIDTH_18_35_2": value  <=  2;
            "WIDTH_18_36_0": value  <=  20;
            "WIDTH_18_36_1": value  <=  20;
            "WIDTH_18_37_0": value  <=  8;
            "WIDTH_18_37_1": value  <=  4;
            "WIDTH_18_37_2": value  <=  4;
            "WIDTH_18_38_0": value  <=  10;
            "WIDTH_18_38_1": value  <=  10;
            "WIDTH_18_39_0": value  <=  2;
            "WIDTH_18_39_1": value  <=  1;
            "WIDTH_18_39_2": value  <=  1;
            "WIDTH_18_40_0": value  <=  2;
            "WIDTH_18_40_1": value  <=  1;
            "WIDTH_18_40_2": value  <=  1;
            "WIDTH_18_41_0": value  <=  3;
            "WIDTH_18_41_1": value  <=  3;
            "WIDTH_18_42_0": value  <=  6;
            "WIDTH_18_42_1": value  <=  2;
            "WIDTH_18_43_0": value  <=  20;
            "WIDTH_18_43_1": value  <=  20;
            "WIDTH_18_44_0": value  <=  8;
            "WIDTH_18_44_1": value  <=  4;
            "WIDTH_18_44_2": value  <=  4;
            "WIDTH_18_45_0": value  <=  18;
            "WIDTH_18_45_1": value  <=  6;
            "WIDTH_18_46_0": value  <=  6;
            "WIDTH_18_46_1": value  <=  6;
            "WIDTH_18_47_0": value  <=  3;
            "WIDTH_18_47_1": value  <=  1;
            "WIDTH_18_48_0": value  <=  6;
            "WIDTH_18_48_1": value  <=  2;
            "WIDTH_18_49_0": value  <=  4;
            "WIDTH_18_49_1": value  <=  4;
            "WIDTH_18_50_0": value  <=  18;
            "WIDTH_18_50_1": value  <=  9;
            "WIDTH_18_51_0": value  <=  1;
            "WIDTH_18_51_1": value  <=  1;
            "WIDTH_18_52_0": value  <=  1;
            "WIDTH_18_52_1": value  <=  1;
            "WIDTH_18_53_0": value  <=  1;
            "WIDTH_18_53_1": value  <=  1;
            "WIDTH_18_54_0": value  <=  1;
            "WIDTH_18_54_1": value  <=  1;
            "WIDTH_18_55_0": value  <=  4;
            "WIDTH_18_55_1": value  <=  4;
            "WIDTH_18_56_0": value  <=  7;
            "WIDTH_18_56_1": value  <=  7;
            "WIDTH_18_57_0": value  <=  6;
            "WIDTH_18_57_1": value  <=  3;
            "WIDTH_18_58_0": value  <=  2;
            "WIDTH_18_58_1": value  <=  2;
            "WIDTH_18_59_0": value  <=  2;
            "WIDTH_18_59_1": value  <=  2;
            "WIDTH_18_60_0": value  <=  8;
            "WIDTH_18_60_1": value  <=  8;
            "WIDTH_18_61_0": value  <=  20;
            "WIDTH_18_61_1": value  <=  10;
            "WIDTH_18_61_2": value  <=  10;
            "WIDTH_18_62_0": value  <=  2;
            "WIDTH_18_62_1": value  <=  1;
            "WIDTH_18_63_0": value  <=  15;
            "WIDTH_18_63_1": value  <=  5;
            "WIDTH_18_64_0": value  <=  12;
            "WIDTH_18_64_1": value  <=  6;
            "WIDTH_18_65_0": value  <=  2;
            "WIDTH_18_65_1": value  <=  1;
            "WIDTH_18_66_0": value  <=  2;
            "WIDTH_18_66_1": value  <=  1;
            "WIDTH_18_67_0": value  <=  4;
            "WIDTH_18_67_1": value  <=  2;
            "WIDTH_18_67_2": value  <=  2;
            "WIDTH_18_68_0": value  <=  10;
            "WIDTH_18_68_1": value  <=  10;
            "WIDTH_18_69_0": value  <=  3;
            "WIDTH_18_69_1": value  <=  3;
            "WIDTH_18_70_0": value  <=  4;
            "WIDTH_18_70_1": value  <=  2;
            "WIDTH_18_70_2": value  <=  2;
            "WIDTH_18_71_0": value  <=  2;
            "WIDTH_18_71_1": value  <=  2;
            "WIDTH_18_72_0": value  <=  1;
            "WIDTH_18_72_1": value  <=  1;
            "WIDTH_18_73_0": value  <=  7;
            "WIDTH_18_73_1": value  <=  7;
            "WIDTH_18_74_0": value  <=  2;
            "WIDTH_18_74_1": value  <=  2;
            "WIDTH_18_75_0": value  <=  3;
            "WIDTH_18_75_1": value  <=  1;
            "WIDTH_18_76_0": value  <=  2;
            "WIDTH_18_76_1": value  <=  1;
            "WIDTH_18_77_0": value  <=  18;
            "WIDTH_18_77_1": value  <=  6;
            "WIDTH_18_78_0": value  <=  8;
            "WIDTH_18_78_1": value  <=  4;
            "WIDTH_18_79_0": value  <=  6;
            "WIDTH_18_79_1": value  <=  3;
            "WIDTH_18_80_0": value  <=  6;
            "WIDTH_18_80_1": value  <=  3;
            "WIDTH_18_81_0": value  <=  3;
            "WIDTH_18_81_1": value  <=  1;
            "WIDTH_18_82_0": value  <=  3;
            "WIDTH_18_82_1": value  <=  1;
            "WIDTH_18_83_0": value  <=  3;
            "WIDTH_18_83_1": value  <=  1;
            "WIDTH_18_84_0": value  <=  3;
            "WIDTH_18_84_1": value  <=  3;
            "WIDTH_18_85_0": value  <=  3;
            "WIDTH_18_85_1": value  <=  1;
            "WIDTH_18_86_0": value  <=  18;
            "WIDTH_18_86_1": value  <=  18;
            "WIDTH_18_87_0": value  <=  3;
            "WIDTH_18_87_1": value  <=  1;
            "WIDTH_18_88_0": value  <=  2;
            "WIDTH_18_88_1": value  <=  2;
            "WIDTH_18_89_0": value  <=  3;
            "WIDTH_18_89_1": value  <=  1;
            "WIDTH_18_90_0": value  <=  3;
            "WIDTH_18_90_1": value  <=  1;
            "WIDTH_18_91_0": value  <=  3;
            "WIDTH_18_91_1": value  <=  1;
            "WIDTH_18_92_0": value  <=  1;
            "WIDTH_18_92_1": value  <=  1;
            "WIDTH_18_93_0": value  <=  2;
            "WIDTH_18_93_1": value  <=  1;
            "WIDTH_18_94_0": value  <=  2;
            "WIDTH_18_94_1": value  <=  1;
            "WIDTH_18_95_0": value  <=  3;
            "WIDTH_18_95_1": value  <=  1;
            "WIDTH_18_96_0": value  <=  3;
            "WIDTH_18_96_1": value  <=  1;
            "WIDTH_18_97_0": value  <=  2;
            "WIDTH_18_97_1": value  <=  1;
            "WIDTH_18_97_2": value  <=  1;
            "WIDTH_18_98_0": value  <=  2;
            "WIDTH_18_98_1": value  <=  1;
            "WIDTH_18_98_2": value  <=  1;
            "WIDTH_18_99_0": value  <=  3;
            "WIDTH_18_99_1": value  <=  1;
            "WIDTH_18_100_0": value  <=  3;
            "WIDTH_18_100_1": value  <=  1;
            "WIDTH_18_101_0": value  <=  6;
            "WIDTH_18_101_1": value  <=  2;
            "WIDTH_18_102_0": value  <=  6;
            "WIDTH_18_102_1": value  <=  2;
            "WIDTH_18_103_0": value  <=  16;
            "WIDTH_18_103_1": value  <=  8;
            "WIDTH_18_103_2": value  <=  8;
            "WIDTH_18_104_0": value  <=  5;
            "WIDTH_18_104_1": value  <=  5;
            "WIDTH_18_105_0": value  <=  3;
            "WIDTH_18_105_1": value  <=  1;
            "WIDTH_18_106_0": value  <=  4;
            "WIDTH_18_106_1": value  <=  4;
            "WIDTH_18_107_0": value  <=  2;
            "WIDTH_18_107_1": value  <=  1;
            "WIDTH_18_108_0": value  <=  15;
            "WIDTH_18_108_1": value  <=  5;
            "WIDTH_18_109_0": value  <=  7;
            "WIDTH_18_109_1": value  <=  7;
            "WIDTH_18_110_0": value  <=  16;
            "WIDTH_18_110_1": value  <=  8;
            "WIDTH_18_110_2": value  <=  8;
            "WIDTH_18_111_0": value  <=  8;
            "WIDTH_18_111_1": value  <=  8;
            "WIDTH_18_112_0": value  <=  3;
            "WIDTH_18_112_1": value  <=  3;
            "WIDTH_18_113_0": value  <=  14;
            "WIDTH_18_113_1": value  <=  7;
            "WIDTH_18_113_2": value  <=  7;
            "WIDTH_18_114_0": value  <=  3;
            "WIDTH_18_114_1": value  <=  3;
            "WIDTH_18_115_0": value  <=  6;
            "WIDTH_18_115_1": value  <=  2;
            "WIDTH_18_116_0": value  <=  7;
            "WIDTH_18_116_1": value  <=  7;
            "WIDTH_18_117_0": value  <=  6;
            "WIDTH_18_117_1": value  <=  6;
            "WIDTH_18_118_0": value  <=  2;
            "WIDTH_18_118_1": value  <=  2;
            "WIDTH_18_119_0": value  <=  20;
            "WIDTH_18_119_1": value  <=  20;
            "WIDTH_18_120_0": value  <=  6;
            "WIDTH_18_120_1": value  <=  2;
            "WIDTH_18_121_0": value  <=  6;
            "WIDTH_18_121_1": value  <=  2;
            "WIDTH_18_122_0": value  <=  6;
            "WIDTH_18_122_1": value  <=  2;
            "WIDTH_18_123_0": value  <=  3;
            "WIDTH_18_123_1": value  <=  1;
            "WIDTH_18_124_0": value  <=  3;
            "WIDTH_18_124_1": value  <=  1;
            "WIDTH_18_125_0": value  <=  16;
            "WIDTH_18_125_1": value  <=  16;
            "WIDTH_18_126_0": value  <=  15;
            "WIDTH_18_126_1": value  <=  15;
            "WIDTH_18_127_0": value  <=  5;
            "WIDTH_18_127_1": value  <=  5;
            "WIDTH_18_128_0": value  <=  2;
            "WIDTH_18_128_1": value  <=  1;
            "WIDTH_18_129_0": value  <=  9;
            "WIDTH_18_129_1": value  <=  9;
            "WIDTH_18_130_0": value  <=  15;
            "WIDTH_18_130_1": value  <=  5;
            "WIDTH_18_131_0": value  <=  3;
            "WIDTH_18_131_1": value  <=  1;
            "WIDTH_18_132_0": value  <=  20;
            "WIDTH_18_132_1": value  <=  20;
            "WIDTH_18_133_0": value  <=  3;
            "WIDTH_18_133_1": value  <=  1;
            "WIDTH_18_134_0": value  <=  3;
            "WIDTH_18_134_1": value  <=  1;
            "WIDTH_18_135_0": value  <=  3;
            "WIDTH_18_135_1": value  <=  3;
            "WIDTH_18_136_0": value  <=  4;
            "WIDTH_18_136_1": value  <=  4;
            "WIDTH_18_137_0": value  <=  2;
            "WIDTH_18_137_1": value  <=  2;
            "WIDTH_18_138_0": value  <=  4;
            "WIDTH_18_138_1": value  <=  4;
            "WIDTH_18_139_0": value  <=  8;
            "WIDTH_18_139_1": value  <=  4;
            "WIDTH_18_139_2": value  <=  4;
            "WIDTH_18_140_0": value  <=  8;
            "WIDTH_18_140_1": value  <=  8;
            "WIDTH_18_141_0": value  <=  6;
            "WIDTH_18_141_1": value  <=  2;
            "WIDTH_18_142_0": value  <=  2;
            "WIDTH_18_142_1": value  <=  2;
            "WIDTH_18_143_0": value  <=  2;
            "WIDTH_18_143_1": value  <=  1;
            "WIDTH_18_144_0": value  <=  6;
            "WIDTH_18_144_1": value  <=  2;
            "WIDTH_18_145_0": value  <=  14;
            "WIDTH_18_145_1": value  <=  7;
            "WIDTH_18_145_2": value  <=  7;
            "WIDTH_18_146_0": value  <=  4;
            "WIDTH_18_146_1": value  <=  2;
            "WIDTH_18_146_2": value  <=  2;
            "WIDTH_18_147_0": value  <=  3;
            "WIDTH_18_147_1": value  <=  3;
            "WIDTH_18_148_0": value  <=  10;
            "WIDTH_18_148_1": value  <=  5;
            "WIDTH_18_148_2": value  <=  5;
            "WIDTH_18_149_0": value  <=  2;
            "WIDTH_18_149_1": value  <=  2;
            "WIDTH_18_150_0": value  <=  2;
            "WIDTH_18_150_1": value  <=  2;
            "WIDTH_18_151_0": value  <=  4;
            "WIDTH_18_151_1": value  <=  2;
            "WIDTH_18_151_2": value  <=  2;
            "WIDTH_18_152_0": value  <=  7;
            "WIDTH_18_152_1": value  <=  7;
            "WIDTH_18_153_0": value  <=  18;
            "WIDTH_18_153_1": value  <=  9;
            "WIDTH_18_153_2": value  <=  9;
            "WIDTH_18_154_0": value  <=  18;
            "WIDTH_18_154_1": value  <=  9;
            "WIDTH_18_154_2": value  <=  9;
            "WIDTH_18_155_0": value  <=  4;
            "WIDTH_18_155_1": value  <=  2;
            "WIDTH_18_155_2": value  <=  2;
            "WIDTH_18_156_0": value  <=  4;
            "WIDTH_18_156_1": value  <=  2;
            "WIDTH_18_156_2": value  <=  2;
            "WIDTH_18_157_0": value  <=  2;
            "WIDTH_18_157_1": value  <=  2;
            "WIDTH_18_158_0": value  <=  10;
            "WIDTH_18_158_1": value  <=  5;
            "WIDTH_18_158_2": value  <=  5;
            "WIDTH_18_159_0": value  <=  4;
            "WIDTH_18_159_1": value  <=  2;
            "WIDTH_18_159_2": value  <=  2;
            "WIDTH_18_160_0": value  <=  6;
            "WIDTH_18_160_1": value  <=  3;
            "WIDTH_18_161_0": value  <=  4;
            "WIDTH_18_161_1": value  <=  2;
            "WIDTH_18_161_2": value  <=  2;
            "WIDTH_18_162_0": value  <=  2;
            "WIDTH_18_162_1": value  <=  1;
            "WIDTH_18_163_0": value  <=  1;
            "WIDTH_18_163_1": value  <=  1;
            "WIDTH_18_164_0": value  <=  6;
            "WIDTH_18_164_1": value  <=  3;
            "WIDTH_18_165_0": value  <=  4;
            "WIDTH_18_165_1": value  <=  2;
            "WIDTH_18_165_2": value  <=  2;
            "WIDTH_18_166_0": value  <=  4;
            "WIDTH_18_166_1": value  <=  2;
            "WIDTH_18_166_2": value  <=  2;
            "WIDTH_18_167_0": value  <=  4;
            "WIDTH_18_167_1": value  <=  2;
            "WIDTH_18_167_2": value  <=  2;
            "WIDTH_18_168_0": value  <=  6;
            "WIDTH_18_168_1": value  <=  6;
            "WIDTH_18_169_0": value  <=  4;
            "WIDTH_18_169_1": value  <=  2;
            "WIDTH_18_169_2": value  <=  2;
            "WIDTH_18_170_0": value  <=  3;
            "WIDTH_18_170_1": value  <=  1;
            "WIDTH_18_171_0": value  <=  4;
            "WIDTH_18_171_1": value  <=  2;
            "WIDTH_18_171_2": value  <=  2;
            "WIDTH_18_172_0": value  <=  4;
            "WIDTH_18_172_1": value  <=  2;
            "WIDTH_18_172_2": value  <=  2;
            "WIDTH_18_173_0": value  <=  2;
            "WIDTH_18_173_1": value  <=  1;
            "WIDTH_18_173_2": value  <=  1;
            "WIDTH_18_174_0": value  <=  3;
            "WIDTH_18_174_1": value  <=  1;
            "WIDTH_18_175_0": value  <=  17;
            "WIDTH_18_175_1": value  <=  17;
            "WIDTH_18_176_0": value  <=  20;
            "WIDTH_18_176_1": value  <=  20;
            "WIDTH_19_0_0": value  <=  8;
            "WIDTH_19_0_1": value  <=  4;
            "WIDTH_19_1_0": value  <=  4;
            "WIDTH_19_1_1": value  <=  4;
            "WIDTH_19_2_0": value  <=  6;
            "WIDTH_19_2_1": value  <=  3;
            "WIDTH_19_2_2": value  <=  3;
            "WIDTH_19_3_0": value  <=  4;
            "WIDTH_19_3_1": value  <=  4;
            "WIDTH_19_4_0": value  <=  1;
            "WIDTH_19_4_1": value  <=  1;
            "WIDTH_19_5_0": value  <=  12;
            "WIDTH_19_5_1": value  <=  4;
            "WIDTH_19_6_0": value  <=  4;
            "WIDTH_19_6_1": value  <=  2;
            "WIDTH_19_6_2": value  <=  2;
            "WIDTH_19_7_0": value  <=  17;
            "WIDTH_19_7_1": value  <=  17;
            "WIDTH_19_8_0": value  <=  16;
            "WIDTH_19_8_1": value  <=  16;
            "WIDTH_19_9_0": value  <=  5;
            "WIDTH_19_9_1": value  <=  5;
            "WIDTH_19_10_0": value  <=  2;
            "WIDTH_19_10_1": value  <=  1;
            "WIDTH_19_11_0": value  <=  16;
            "WIDTH_19_11_1": value  <=  16;
            "WIDTH_19_12_0": value  <=  5;
            "WIDTH_19_12_1": value  <=  5;
            "WIDTH_19_13_0": value  <=  3;
            "WIDTH_19_13_1": value  <=  1;
            "WIDTH_19_14_0": value  <=  3;
            "WIDTH_19_14_1": value  <=  1;
            "WIDTH_19_15_0": value  <=  3;
            "WIDTH_19_15_1": value  <=  3;
            "WIDTH_19_16_0": value  <=  5;
            "WIDTH_19_16_1": value  <=  5;
            "WIDTH_19_17_0": value  <=  4;
            "WIDTH_19_17_1": value  <=  4;
            "WIDTH_19_18_0": value  <=  12;
            "WIDTH_19_18_1": value  <=  4;
            "WIDTH_19_19_0": value  <=  6;
            "WIDTH_19_19_1": value  <=  6;
            "WIDTH_19_20_0": value  <=  8;
            "WIDTH_19_20_1": value  <=  4;
            "WIDTH_19_20_2": value  <=  4;
            "WIDTH_19_21_0": value  <=  3;
            "WIDTH_19_21_1": value  <=  1;
            "WIDTH_19_22_0": value  <=  3;
            "WIDTH_19_22_1": value  <=  1;
            "WIDTH_19_23_0": value  <=  3;
            "WIDTH_19_23_1": value  <=  3;
            "WIDTH_19_24_0": value  <=  6;
            "WIDTH_19_24_1": value  <=  6;
            "WIDTH_19_25_0": value  <=  3;
            "WIDTH_19_25_1": value  <=  3;
            "WIDTH_19_26_0": value  <=  2;
            "WIDTH_19_26_1": value  <=  2;
            "WIDTH_19_27_0": value  <=  6;
            "WIDTH_19_27_1": value  <=  6;
            "WIDTH_19_28_0": value  <=  3;
            "WIDTH_19_28_1": value  <=  3;
            "WIDTH_19_29_0": value  <=  3;
            "WIDTH_19_29_1": value  <=  1;
            "WIDTH_19_30_0": value  <=  2;
            "WIDTH_19_30_1": value  <=  2;
            "WIDTH_19_31_0": value  <=  3;
            "WIDTH_19_31_1": value  <=  3;
            "WIDTH_19_32_0": value  <=  2;
            "WIDTH_19_32_1": value  <=  2;
            "WIDTH_19_33_0": value  <=  6;
            "WIDTH_19_33_1": value  <=  6;
            "WIDTH_19_34_0": value  <=  16;
            "WIDTH_19_34_1": value  <=  16;
            "WIDTH_19_35_0": value  <=  6;
            "WIDTH_19_35_1": value  <=  6;
            "WIDTH_19_36_0": value  <=  5;
            "WIDTH_19_36_1": value  <=  5;
            "WIDTH_19_37_0": value  <=  4;
            "WIDTH_19_37_1": value  <=  4;
            "WIDTH_19_38_0": value  <=  3;
            "WIDTH_19_38_1": value  <=  3;
            "WIDTH_19_39_0": value  <=  4;
            "WIDTH_19_39_1": value  <=  4;
            "WIDTH_19_40_0": value  <=  1;
            "WIDTH_19_40_1": value  <=  1;
            "WIDTH_19_41_0": value  <=  4;
            "WIDTH_19_41_1": value  <=  4;
            "WIDTH_19_42_0": value  <=  8;
            "WIDTH_19_42_1": value  <=  8;
            "WIDTH_19_43_0": value  <=  4;
            "WIDTH_19_43_1": value  <=  4;
            "WIDTH_19_44_0": value  <=  9;
            "WIDTH_19_44_1": value  <=  3;
            "WIDTH_19_45_0": value  <=  4;
            "WIDTH_19_45_1": value  <=  4;
            "WIDTH_19_46_0": value  <=  4;
            "WIDTH_19_46_1": value  <=  4;
            "WIDTH_19_47_0": value  <=  9;
            "WIDTH_19_47_1": value  <=  3;
            "WIDTH_19_48_0": value  <=  1;
            "WIDTH_19_48_1": value  <=  1;
            "WIDTH_19_49_0": value  <=  6;
            "WIDTH_19_49_1": value  <=  3;
            "WIDTH_19_50_0": value  <=  3;
            "WIDTH_19_50_1": value  <=  1;
            "WIDTH_19_51_0": value  <=  3;
            "WIDTH_19_51_1": value  <=  1;
            "WIDTH_19_52_0": value  <=  3;
            "WIDTH_19_52_1": value  <=  1;
            "WIDTH_19_53_0": value  <=  11;
            "WIDTH_19_53_1": value  <=  11;
            "WIDTH_19_54_0": value  <=  10;
            "WIDTH_19_54_1": value  <=  5;
            "WIDTH_19_55_0": value  <=  3;
            "WIDTH_19_55_1": value  <=  1;
            "WIDTH_19_56_0": value  <=  3;
            "WIDTH_19_56_1": value  <=  1;
            "WIDTH_19_57_0": value  <=  4;
            "WIDTH_19_57_1": value  <=  2;
            "WIDTH_19_58_0": value  <=  4;
            "WIDTH_19_58_1": value  <=  2;
            "WIDTH_19_59_0": value  <=  2;
            "WIDTH_19_59_1": value  <=  2;
            "WIDTH_19_60_0": value  <=  3;
            "WIDTH_19_60_1": value  <=  1;
            "WIDTH_19_61_0": value  <=  6;
            "WIDTH_19_61_1": value  <=  6;
            "WIDTH_19_62_0": value  <=  12;
            "WIDTH_19_62_1": value  <=  6;
            "WIDTH_19_62_2": value  <=  6;
            "WIDTH_19_63_0": value  <=  8;
            "WIDTH_19_63_1": value  <=  4;
            "WIDTH_19_63_2": value  <=  4;
            "WIDTH_19_64_0": value  <=  15;
            "WIDTH_19_64_1": value  <=  5;
            "WIDTH_19_65_0": value  <=  4;
            "WIDTH_19_65_1": value  <=  2;
            "WIDTH_19_66_0": value  <=  2;
            "WIDTH_19_66_1": value  <=  2;
            "WIDTH_19_67_0": value  <=  4;
            "WIDTH_19_67_1": value  <=  4;
            "WIDTH_19_68_0": value  <=  2;
            "WIDTH_19_68_1": value  <=  2;
            "WIDTH_19_69_0": value  <=  2;
            "WIDTH_19_69_1": value  <=  2;
            "WIDTH_19_70_0": value  <=  4;
            "WIDTH_19_70_1": value  <=  2;
            "WIDTH_19_70_2": value  <=  2;
            "WIDTH_19_71_0": value  <=  2;
            "WIDTH_19_71_1": value  <=  1;
            "WIDTH_19_71_2": value  <=  1;
            "WIDTH_19_72_0": value  <=  3;
            "WIDTH_19_72_1": value  <=  1;
            "WIDTH_19_73_0": value  <=  2;
            "WIDTH_19_73_1": value  <=  1;
            "WIDTH_19_73_2": value  <=  1;
            "WIDTH_19_74_0": value  <=  6;
            "WIDTH_19_74_1": value  <=  6;
            "WIDTH_19_75_0": value  <=  2;
            "WIDTH_19_75_1": value  <=  1;
            "WIDTH_19_75_2": value  <=  1;
            "WIDTH_19_76_0": value  <=  2;
            "WIDTH_19_76_1": value  <=  1;
            "WIDTH_19_76_2": value  <=  1;
            "WIDTH_19_77_0": value  <=  8;
            "WIDTH_19_77_1": value  <=  4;
            "WIDTH_19_78_0": value  <=  8;
            "WIDTH_19_78_1": value  <=  4;
            "WIDTH_19_79_0": value  <=  4;
            "WIDTH_19_79_1": value  <=  2;
            "WIDTH_19_80_0": value  <=  4;
            "WIDTH_19_80_1": value  <=  2;
            "WIDTH_19_81_0": value  <=  4;
            "WIDTH_19_81_1": value  <=  2;
            "WIDTH_19_81_2": value  <=  2;
            "WIDTH_19_82_0": value  <=  3;
            "WIDTH_19_82_1": value  <=  1;
            "WIDTH_19_83_0": value  <=  4;
            "WIDTH_19_83_1": value  <=  2;
            "WIDTH_19_83_2": value  <=  2;
            "WIDTH_19_84_0": value  <=  2;
            "WIDTH_19_84_1": value  <=  2;
            "WIDTH_19_85_0": value  <=  15;
            "WIDTH_19_85_1": value  <=  15;
            "WIDTH_19_86_0": value  <=  2;
            "WIDTH_19_86_1": value  <=  1;
            "WIDTH_19_86_2": value  <=  1;
            "WIDTH_19_87_0": value  <=  2;
            "WIDTH_19_87_1": value  <=  2;
            "WIDTH_19_88_0": value  <=  3;
            "WIDTH_19_88_1": value  <=  1;
            "WIDTH_19_89_0": value  <=  3;
            "WIDTH_19_89_1": value  <=  1;
            "WIDTH_19_90_0": value  <=  3;
            "WIDTH_19_90_1": value  <=  1;
            "WIDTH_19_91_0": value  <=  4;
            "WIDTH_19_91_1": value  <=  2;
            "WIDTH_19_91_2": value  <=  2;
            "WIDTH_19_92_0": value  <=  2;
            "WIDTH_19_92_1": value  <=  2;
            "WIDTH_19_93_0": value  <=  18;
            "WIDTH_19_93_1": value  <=  6;
            "WIDTH_19_94_0": value  <=  4;
            "WIDTH_19_94_1": value  <=  2;
            "WIDTH_19_95_0": value  <=  12;
            "WIDTH_19_95_1": value  <=  6;
            "WIDTH_19_96_0": value  <=  18;
            "WIDTH_19_96_1": value  <=  6;
            "WIDTH_19_97_0": value  <=  2;
            "WIDTH_19_97_1": value  <=  2;
            "WIDTH_19_98_0": value  <=  1;
            "WIDTH_19_98_1": value  <=  1;
            "WIDTH_19_99_0": value  <=  2;
            "WIDTH_19_99_1": value  <=  2;
            "WIDTH_19_100_0": value  <=  2;
            "WIDTH_19_100_1": value  <=  2;
            "WIDTH_19_101_0": value  <=  3;
            "WIDTH_19_101_1": value  <=  3;
            "WIDTH_19_102_0": value  <=  4;
            "WIDTH_19_102_1": value  <=  2;
            "WIDTH_19_103_0": value  <=  6;
            "WIDTH_19_103_1": value  <=  3;
            "WIDTH_19_103_2": value  <=  3;
            "WIDTH_19_104_0": value  <=  12;
            "WIDTH_19_104_1": value  <=  12;
            "WIDTH_19_105_0": value  <=  4;
            "WIDTH_19_105_1": value  <=  2;
            "WIDTH_19_105_2": value  <=  2;
            "WIDTH_19_106_0": value  <=  10;
            "WIDTH_19_106_1": value  <=  5;
            "WIDTH_19_106_2": value  <=  5;
            "WIDTH_19_107_0": value  <=  4;
            "WIDTH_19_107_1": value  <=  4;
            "WIDTH_19_108_0": value  <=  8;
            "WIDTH_19_108_1": value  <=  8;
            "WIDTH_19_109_0": value  <=  5;
            "WIDTH_19_109_1": value  <=  5;
            "WIDTH_19_110_0": value  <=  4;
            "WIDTH_19_110_1": value  <=  4;
            "WIDTH_19_111_0": value  <=  6;
            "WIDTH_19_111_1": value  <=  6;
            "WIDTH_19_112_0": value  <=  8;
            "WIDTH_19_112_1": value  <=  4;
            "WIDTH_19_112_2": value  <=  4;
            "WIDTH_19_113_0": value  <=  3;
            "WIDTH_19_113_1": value  <=  3;
            "WIDTH_19_114_0": value  <=  4;
            "WIDTH_19_114_1": value  <=  4;
            "WIDTH_19_115_0": value  <=  6;
            "WIDTH_19_115_1": value  <=  6;
            "WIDTH_19_116_0": value  <=  3;
            "WIDTH_19_116_1": value  <=  1;
            "WIDTH_19_117_0": value  <=  3;
            "WIDTH_19_117_1": value  <=  3;
            "WIDTH_19_118_0": value  <=  6;
            "WIDTH_19_118_1": value  <=  6;
            "WIDTH_19_119_0": value  <=  3;
            "WIDTH_19_119_1": value  <=  1;
            "WIDTH_19_120_0": value  <=  3;
            "WIDTH_19_120_1": value  <=  1;
            "WIDTH_19_121_0": value  <=  1;
            "WIDTH_19_121_1": value  <=  1;
            "WIDTH_19_122_0": value  <=  4;
            "WIDTH_19_122_1": value  <=  2;
            "WIDTH_19_123_0": value  <=  3;
            "WIDTH_19_123_1": value  <=  3;
            "WIDTH_19_124_0": value  <=  3;
            "WIDTH_19_124_1": value  <=  3;
            "WIDTH_19_125_0": value  <=  6;
            "WIDTH_19_125_1": value  <=  3;
            "WIDTH_19_125_2": value  <=  3;
            "WIDTH_19_126_0": value  <=  6;
            "WIDTH_19_126_1": value  <=  3;
            "WIDTH_19_126_2": value  <=  3;
            "WIDTH_19_127_0": value  <=  4;
            "WIDTH_19_127_1": value  <=  4;
            "WIDTH_19_128_0": value  <=  6;
            "WIDTH_19_128_1": value  <=  2;
            "WIDTH_19_129_0": value  <=  3;
            "WIDTH_19_129_1": value  <=  1;
            "WIDTH_19_130_0": value  <=  3;
            "WIDTH_19_130_1": value  <=  1;
            "WIDTH_19_131_0": value  <=  6;
            "WIDTH_19_131_1": value  <=  2;
            "WIDTH_19_132_0": value  <=  8;
            "WIDTH_19_132_1": value  <=  4;
            "WIDTH_19_133_0": value  <=  2;
            "WIDTH_19_133_1": value  <=  1;
            "WIDTH_19_134_0": value  <=  3;
            "WIDTH_19_134_1": value  <=  1;
            "WIDTH_19_135_0": value  <=  6;
            "WIDTH_19_135_1": value  <=  2;
            "WIDTH_19_136_0": value  <=  3;
            "WIDTH_19_136_1": value  <=  1;
            "WIDTH_19_137_0": value  <=  3;
            "WIDTH_19_137_1": value  <=  1;
            "WIDTH_19_138_0": value  <=  6;
            "WIDTH_19_138_1": value  <=  2;
            "WIDTH_19_139_0": value  <=  3;
            "WIDTH_19_139_1": value  <=  3;
            "WIDTH_19_140_0": value  <=  4;
            "WIDTH_19_140_1": value  <=  4;
            "WIDTH_19_141_0": value  <=  3;
            "WIDTH_19_141_1": value  <=  3;
            "WIDTH_19_142_0": value  <=  3;
            "WIDTH_19_142_1": value  <=  3;
            "WIDTH_19_143_0": value  <=  6;
            "WIDTH_19_143_1": value  <=  3;
            "WIDTH_19_143_2": value  <=  3;
            "WIDTH_19_144_0": value  <=  5;
            "WIDTH_19_144_1": value  <=  5;
            "WIDTH_19_145_0": value  <=  2;
            "WIDTH_19_145_1": value  <=  1;
            "WIDTH_19_145_2": value  <=  1;
            "WIDTH_19_146_0": value  <=  3;
            "WIDTH_19_146_1": value  <=  3;
            "WIDTH_19_147_0": value  <=  3;
            "WIDTH_19_147_1": value  <=  3;
            "WIDTH_19_148_0": value  <=  3;
            "WIDTH_19_148_1": value  <=  3;
            "WIDTH_19_149_0": value  <=  9;
            "WIDTH_19_149_1": value  <=  9;
            "WIDTH_19_150_0": value  <=  3;
            "WIDTH_19_150_1": value  <=  1;
            "WIDTH_19_151_0": value  <=  12;
            "WIDTH_19_151_1": value  <=  4;
            "WIDTH_19_152_0": value  <=  2;
            "WIDTH_19_152_1": value  <=  1;
            "WIDTH_19_152_2": value  <=  1;
            "WIDTH_19_153_0": value  <=  3;
            "WIDTH_19_153_1": value  <=  3;
            "WIDTH_19_154_0": value  <=  3;
            "WIDTH_19_154_1": value  <=  3;
            "WIDTH_19_155_0": value  <=  6;
            "WIDTH_19_155_1": value  <=  3;
            "WIDTH_19_155_2": value  <=  3;
            "WIDTH_19_156_0": value  <=  15;
            "WIDTH_19_156_1": value  <=  5;
            "WIDTH_19_157_0": value  <=  18;
            "WIDTH_19_157_1": value  <=  6;
            "WIDTH_19_158_0": value  <=  4;
            "WIDTH_19_158_1": value  <=  2;
            "WIDTH_19_159_0": value  <=  12;
            "WIDTH_19_159_1": value  <=  4;
            "WIDTH_19_160_0": value  <=  12;
            "WIDTH_19_160_1": value  <=  4;
            "WIDTH_19_161_0": value  <=  12;
            "WIDTH_19_161_1": value  <=  6;
            "WIDTH_19_161_2": value  <=  6;
            "WIDTH_19_162_0": value  <=  6;
            "WIDTH_19_162_1": value  <=  3;
            "WIDTH_19_162_2": value  <=  3;
            "WIDTH_19_163_0": value  <=  2;
            "WIDTH_19_163_1": value  <=  2;
            "WIDTH_19_164_0": value  <=  20;
            "WIDTH_19_164_1": value  <=  10;
            "WIDTH_19_164_2": value  <=  10;
            "WIDTH_19_165_0": value  <=  12;
            "WIDTH_19_165_1": value  <=  6;
            "WIDTH_19_165_2": value  <=  6;
            "WIDTH_19_166_0": value  <=  3;
            "WIDTH_19_166_1": value  <=  3;
            "WIDTH_19_167_0": value  <=  2;
            "WIDTH_19_167_1": value  <=  2;
            "WIDTH_19_168_0": value  <=  2;
            "WIDTH_19_168_1": value  <=  1;
            "WIDTH_19_168_2": value  <=  1;
            "WIDTH_19_169_0": value  <=  14;
            "WIDTH_19_169_1": value  <=  7;
            "WIDTH_19_169_2": value  <=  7;
            "WIDTH_19_170_0": value  <=  4;
            "WIDTH_19_170_1": value  <=  4;
            "WIDTH_19_171_0": value  <=  6;
            "WIDTH_19_171_1": value  <=  2;
            "WIDTH_19_172_0": value  <=  1;
            "WIDTH_19_172_1": value  <=  1;
            "WIDTH_19_173_0": value  <=  6;
            "WIDTH_19_173_1": value  <=  3;
            "WIDTH_19_173_2": value  <=  3;
            "WIDTH_19_174_0": value  <=  6;
            "WIDTH_19_174_1": value  <=  3;
            "WIDTH_19_174_2": value  <=  3;
            "WIDTH_19_175_0": value  <=  6;
            "WIDTH_19_175_1": value  <=  2;
            "WIDTH_19_176_0": value  <=  8;
            "WIDTH_19_176_1": value  <=  4;
            "WIDTH_19_176_2": value  <=  4;
            "WIDTH_19_177_0": value  <=  8;
            "WIDTH_19_177_1": value  <=  4;
            "WIDTH_19_177_2": value  <=  4;
            "WIDTH_19_178_0": value  <=  6;
            "WIDTH_19_178_1": value  <=  2;
            "WIDTH_19_179_0": value  <=  4;
            "WIDTH_19_179_1": value  <=  2;
            "WIDTH_19_180_0": value  <=  4;
            "WIDTH_19_180_1": value  <=  2;
            "WIDTH_19_181_0": value  <=  2;
            "WIDTH_19_181_1": value  <=  1;
            "WIDTH_20_0_0": value  <=  4;
            "WIDTH_20_0_1": value  <=  2;
            "WIDTH_20_1_0": value  <=  6;
            "WIDTH_20_1_1": value  <=  2;
            "WIDTH_20_2_0": value  <=  2;
            "WIDTH_20_2_1": value  <=  2;
            "WIDTH_20_3_0": value  <=  2;
            "WIDTH_20_3_1": value  <=  2;
            "WIDTH_20_4_0": value  <=  5;
            "WIDTH_20_4_1": value  <=  5;
            "WIDTH_20_5_0": value  <=  2;
            "WIDTH_20_5_1": value  <=  2;
            "WIDTH_20_6_0": value  <=  2;
            "WIDTH_20_6_1": value  <=  2;
            "WIDTH_20_7_0": value  <=  10;
            "WIDTH_20_7_1": value  <=  5;
            "WIDTH_20_7_2": value  <=  5;
            "WIDTH_20_8_0": value  <=  2;
            "WIDTH_20_8_1": value  <=  1;
            "WIDTH_20_9_0": value  <=  6;
            "WIDTH_20_9_1": value  <=  6;
            "WIDTH_20_10_0": value  <=  16;
            "WIDTH_20_10_1": value  <=  16;
            "WIDTH_20_11_0": value  <=  6;
            "WIDTH_20_11_1": value  <=  6;
            "WIDTH_20_12_0": value  <=  10;
            "WIDTH_20_12_1": value  <=  10;
            "WIDTH_20_13_0": value  <=  6;
            "WIDTH_20_13_1": value  <=  6;
            "WIDTH_20_14_0": value  <=  6;
            "WIDTH_20_14_1": value  <=  6;
            "WIDTH_20_15_0": value  <=  4;
            "WIDTH_20_15_1": value  <=  2;
            "WIDTH_20_16_0": value  <=  9;
            "WIDTH_20_16_1": value  <=  9;
            "WIDTH_20_17_0": value  <=  3;
            "WIDTH_20_17_1": value  <=  3;
            "WIDTH_20_18_0": value  <=  6;
            "WIDTH_20_18_1": value  <=  2;
            "WIDTH_20_19_0": value  <=  1;
            "WIDTH_20_19_1": value  <=  1;
            "WIDTH_20_20_0": value  <=  2;
            "WIDTH_20_20_1": value  <=  2;
            "WIDTH_20_21_0": value  <=  2;
            "WIDTH_20_21_1": value  <=  2;
            "WIDTH_20_22_0": value  <=  4;
            "WIDTH_20_22_1": value  <=  2;
            "WIDTH_20_23_0": value  <=  4;
            "WIDTH_20_23_1": value  <=  2;
            "WIDTH_20_24_0": value  <=  20;
            "WIDTH_20_24_1": value  <=  10;
            "WIDTH_20_25_0": value  <=  1;
            "WIDTH_20_25_1": value  <=  1;
            "WIDTH_20_26_0": value  <=  3;
            "WIDTH_20_26_1": value  <=  1;
            "WIDTH_20_27_0": value  <=  3;
            "WIDTH_20_27_1": value  <=  3;
            "WIDTH_20_28_0": value  <=  3;
            "WIDTH_20_28_1": value  <=  3;
            "WIDTH_20_29_0": value  <=  12;
            "WIDTH_20_29_1": value  <=  6;
            "WIDTH_20_29_2": value  <=  6;
            "WIDTH_20_30_0": value  <=  4;
            "WIDTH_20_30_1": value  <=  4;
            "WIDTH_20_31_0": value  <=  14;
            "WIDTH_20_31_1": value  <=  7;
            "WIDTH_20_31_2": value  <=  7;
            "WIDTH_20_32_0": value  <=  2;
            "WIDTH_20_32_1": value  <=  2;
            "WIDTH_20_33_0": value  <=  2;
            "WIDTH_20_33_1": value  <=  2;
            "WIDTH_20_34_0": value  <=  4;
            "WIDTH_20_34_1": value  <=  4;
            "WIDTH_20_35_0": value  <=  1;
            "WIDTH_20_35_1": value  <=  1;
            "WIDTH_20_36_0": value  <=  5;
            "WIDTH_20_36_1": value  <=  5;
            "WIDTH_20_37_0": value  <=  6;
            "WIDTH_20_37_1": value  <=  6;
            "WIDTH_20_38_0": value  <=  4;
            "WIDTH_20_38_1": value  <=  4;
            "WIDTH_20_39_0": value  <=  3;
            "WIDTH_20_39_1": value  <=  1;
            "WIDTH_20_40_0": value  <=  3;
            "WIDTH_20_40_1": value  <=  1;
            "WIDTH_20_41_0": value  <=  3;
            "WIDTH_20_41_1": value  <=  1;
            "WIDTH_20_42_0": value  <=  12;
            "WIDTH_20_42_1": value  <=  4;
            "WIDTH_20_43_0": value  <=  3;
            "WIDTH_20_43_1": value  <=  1;
            "WIDTH_20_44_0": value  <=  2;
            "WIDTH_20_44_1": value  <=  2;
            "WIDTH_20_45_0": value  <=  3;
            "WIDTH_20_45_1": value  <=  1;
            "WIDTH_20_46_0": value  <=  3;
            "WIDTH_20_46_1": value  <=  1;
            "WIDTH_20_47_0": value  <=  18;
            "WIDTH_20_47_1": value  <=  6;
            "WIDTH_20_48_0": value  <=  8;
            "WIDTH_20_48_1": value  <=  4;
            "WIDTH_20_49_0": value  <=  8;
            "WIDTH_20_49_1": value  <=  8;
            "WIDTH_20_50_0": value  <=  8;
            "WIDTH_20_50_1": value  <=  8;
            "WIDTH_20_51_0": value  <=  2;
            "WIDTH_20_51_1": value  <=  2;
            "WIDTH_20_52_0": value  <=  12;
            "WIDTH_20_52_1": value  <=  6;
            "WIDTH_20_52_2": value  <=  6;
            "WIDTH_20_53_0": value  <=  3;
            "WIDTH_20_53_1": value  <=  1;
            "WIDTH_20_54_0": value  <=  3;
            "WIDTH_20_54_1": value  <=  1;
            "WIDTH_20_55_0": value  <=  4;
            "WIDTH_20_55_1": value  <=  2;
            "WIDTH_20_55_2": value  <=  2;
            "WIDTH_20_56_0": value  <=  3;
            "WIDTH_20_56_1": value  <=  1;
            "WIDTH_20_57_0": value  <=  4;
            "WIDTH_20_57_1": value  <=  4;
            "WIDTH_20_58_0": value  <=  3;
            "WIDTH_20_58_1": value  <=  1;
            "WIDTH_20_59_0": value  <=  6;
            "WIDTH_20_59_1": value  <=  6;
            "WIDTH_20_60_0": value  <=  6;
            "WIDTH_20_60_1": value  <=  2;
            "WIDTH_20_61_0": value  <=  2;
            "WIDTH_20_61_1": value  <=  2;
            "WIDTH_20_62_0": value  <=  3;
            "WIDTH_20_62_1": value  <=  1;
            "WIDTH_20_63_0": value  <=  2;
            "WIDTH_20_63_1": value  <=  2;
            "WIDTH_20_64_0": value  <=  4;
            "WIDTH_20_64_1": value  <=  2;
            "WIDTH_20_65_0": value  <=  2;
            "WIDTH_20_65_1": value  <=  2;
            "WIDTH_20_66_0": value  <=  2;
            "WIDTH_20_66_1": value  <=  2;
            "WIDTH_20_67_0": value  <=  2;
            "WIDTH_20_67_1": value  <=  1;
            "WIDTH_20_67_2": value  <=  1;
            "WIDTH_20_68_0": value  <=  2;
            "WIDTH_20_68_1": value  <=  1;
            "WIDTH_20_68_2": value  <=  1;
            "WIDTH_20_69_0": value  <=  3;
            "WIDTH_20_69_1": value  <=  1;
            "WIDTH_20_70_0": value  <=  3;
            "WIDTH_20_70_1": value  <=  1;
            "WIDTH_20_71_0": value  <=  3;
            "WIDTH_20_71_1": value  <=  1;
            "WIDTH_20_72_0": value  <=  2;
            "WIDTH_20_72_1": value  <=  2;
            "WIDTH_20_73_0": value  <=  4;
            "WIDTH_20_73_1": value  <=  4;
            "WIDTH_20_74_0": value  <=  3;
            "WIDTH_20_74_1": value  <=  1;
            "WIDTH_20_75_0": value  <=  8;
            "WIDTH_20_75_1": value  <=  8;
            "WIDTH_20_76_0": value  <=  7;
            "WIDTH_20_76_1": value  <=  7;
            "WIDTH_20_77_0": value  <=  10;
            "WIDTH_20_77_1": value  <=  5;
            "WIDTH_20_77_2": value  <=  5;
            "WIDTH_20_78_0": value  <=  8;
            "WIDTH_20_78_1": value  <=  8;
            "WIDTH_20_79_0": value  <=  4;
            "WIDTH_20_79_1": value  <=  4;
            "WIDTH_20_80_0": value  <=  1;
            "WIDTH_20_80_1": value  <=  1;
            "WIDTH_20_81_0": value  <=  4;
            "WIDTH_20_81_1": value  <=  4;
            "WIDTH_20_82_0": value  <=  4;
            "WIDTH_20_82_1": value  <=  2;
            "WIDTH_20_82_2": value  <=  2;
            "WIDTH_20_83_0": value  <=  4;
            "WIDTH_20_83_1": value  <=  4;
            "WIDTH_20_84_0": value  <=  4;
            "WIDTH_20_84_1": value  <=  4;
            "WIDTH_20_85_0": value  <=  2;
            "WIDTH_20_85_1": value  <=  1;
            "WIDTH_20_86_0": value  <=  6;
            "WIDTH_20_86_1": value  <=  6;
            "WIDTH_20_87_0": value  <=  2;
            "WIDTH_20_87_1": value  <=  1;
            "WIDTH_20_88_0": value  <=  2;
            "WIDTH_20_88_1": value  <=  2;
            "WIDTH_20_89_0": value  <=  3;
            "WIDTH_20_89_1": value  <=  3;
            "WIDTH_20_90_0": value  <=  10;
            "WIDTH_20_90_1": value  <=  5;
            "WIDTH_20_90_2": value  <=  5;
            "WIDTH_20_91_0": value  <=  10;
            "WIDTH_20_91_1": value  <=  5;
            "WIDTH_20_91_2": value  <=  5;
            "WIDTH_20_92_0": value  <=  1;
            "WIDTH_20_92_1": value  <=  1;
            "WIDTH_20_93_0": value  <=  6;
            "WIDTH_20_93_1": value  <=  6;
            "WIDTH_20_94_0": value  <=  3;
            "WIDTH_20_94_1": value  <=  3;
            "WIDTH_20_95_0": value  <=  10;
            "WIDTH_20_95_1": value  <=  10;
            "WIDTH_20_96_0": value  <=  5;
            "WIDTH_20_96_1": value  <=  5;
            "WIDTH_20_97_0": value  <=  3;
            "WIDTH_20_97_1": value  <=  3;
            "WIDTH_20_98_0": value  <=  3;
            "WIDTH_20_98_1": value  <=  3;
            "WIDTH_20_99_0": value  <=  2;
            "WIDTH_20_99_1": value  <=  1;
            "WIDTH_20_100_0": value  <=  6;
            "WIDTH_20_100_1": value  <=  2;
            "WIDTH_20_101_0": value  <=  6;
            "WIDTH_20_101_1": value  <=  3;
            "WIDTH_20_102_0": value  <=  15;
            "WIDTH_20_102_1": value  <=  5;
            "WIDTH_20_103_0": value  <=  8;
            "WIDTH_20_103_1": value  <=  4;
            "WIDTH_20_103_2": value  <=  4;
            "WIDTH_20_104_0": value  <=  3;
            "WIDTH_20_104_1": value  <=  3;
            "WIDTH_20_105_0": value  <=  2;
            "WIDTH_20_105_1": value  <=  2;
            "WIDTH_20_106_0": value  <=  2;
            "WIDTH_20_106_1": value  <=  1;
            "WIDTH_20_107_0": value  <=  7;
            "WIDTH_20_107_1": value  <=  7;
            "WIDTH_20_108_0": value  <=  1;
            "WIDTH_20_108_1": value  <=  1;
            "WIDTH_20_109_0": value  <=  2;
            "WIDTH_20_109_1": value  <=  1;
            "WIDTH_20_109_2": value  <=  1;
            "WIDTH_20_110_0": value  <=  7;
            "WIDTH_20_110_1": value  <=  7;
            "WIDTH_20_111_0": value  <=  2;
            "WIDTH_20_111_1": value  <=  1;
            "WIDTH_20_111_2": value  <=  1;
            "WIDTH_20_112_0": value  <=  8;
            "WIDTH_20_112_1": value  <=  4;
            "WIDTH_20_112_2": value  <=  4;
            "WIDTH_20_113_0": value  <=  8;
            "WIDTH_20_113_1": value  <=  8;
            "WIDTH_20_114_0": value  <=  2;
            "WIDTH_20_114_1": value  <=  2;
            "WIDTH_20_115_0": value  <=  6;
            "WIDTH_20_115_1": value  <=  3;
            "WIDTH_20_115_2": value  <=  3;
            "WIDTH_20_116_0": value  <=  20;
            "WIDTH_20_116_1": value  <=  10;
            "WIDTH_20_116_2": value  <=  10;
            "WIDTH_20_117_0": value  <=  2;
            "WIDTH_20_117_1": value  <=  1;
            "WIDTH_20_117_2": value  <=  1;
            "WIDTH_20_118_0": value  <=  6;
            "WIDTH_20_118_1": value  <=  3;
            "WIDTH_20_119_0": value  <=  6;
            "WIDTH_20_119_1": value  <=  3;
            "WIDTH_20_120_0": value  <=  10;
            "WIDTH_20_120_1": value  <=  5;
            "WIDTH_20_121_0": value  <=  4;
            "WIDTH_20_121_1": value  <=  2;
            "WIDTH_20_122_0": value  <=  2;
            "WIDTH_20_122_1": value  <=  1;
            "WIDTH_20_123_0": value  <=  6;
            "WIDTH_20_123_1": value  <=  3;
            "WIDTH_20_124_0": value  <=  6;
            "WIDTH_20_124_1": value  <=  3;
            "WIDTH_20_125_0": value  <=  18;
            "WIDTH_20_125_1": value  <=  6;
            "WIDTH_20_126_0": value  <=  4;
            "WIDTH_20_126_1": value  <=  2;
            "WIDTH_20_127_0": value  <=  12;
            "WIDTH_20_127_1": value  <=  6;
            "WIDTH_20_127_2": value  <=  6;
            "WIDTH_20_128_0": value  <=  20;
            "WIDTH_20_128_1": value  <=  10;
            "WIDTH_20_128_2": value  <=  10;
            "WIDTH_20_129_0": value  <=  14;
            "WIDTH_20_129_1": value  <=  7;
            "WIDTH_20_129_2": value  <=  7;
            "WIDTH_20_130_0": value  <=  10;
            "WIDTH_20_130_1": value  <=  5;
            "WIDTH_20_130_2": value  <=  5;
            "WIDTH_20_131_0": value  <=  14;
            "WIDTH_20_131_1": value  <=  14;
            "WIDTH_20_132_0": value  <=  2;
            "WIDTH_20_132_1": value  <=  2;
            "WIDTH_20_133_0": value  <=  3;
            "WIDTH_20_133_1": value  <=  1;
            "WIDTH_20_134_0": value  <=  4;
            "WIDTH_20_134_1": value  <=  2;
            "WIDTH_20_134_2": value  <=  2;
            "WIDTH_20_135_0": value  <=  1;
            "WIDTH_20_135_1": value  <=  1;
            "WIDTH_20_136_0": value  <=  4;
            "WIDTH_20_136_1": value  <=  2;
            "WIDTH_20_136_2": value  <=  2;
            "WIDTH_20_137_0": value  <=  8;
            "WIDTH_20_137_1": value  <=  8;
            "WIDTH_20_138_0": value  <=  5;
            "WIDTH_20_138_1": value  <=  5;
            "WIDTH_20_139_0": value  <=  6;
            "WIDTH_20_139_1": value  <=  3;
            "WIDTH_20_139_2": value  <=  3;
            "WIDTH_20_140_0": value  <=  18;
            "WIDTH_20_140_1": value  <=  6;
            "WIDTH_20_141_0": value  <=  6;
            "WIDTH_20_141_1": value  <=  3;
            "WIDTH_20_141_2": value  <=  3;
            "WIDTH_20_142_0": value  <=  1;
            "WIDTH_20_142_1": value  <=  1;
            "WIDTH_20_143_0": value  <=  15;
            "WIDTH_20_143_1": value  <=  15;
            "WIDTH_20_144_0": value  <=  6;
            "WIDTH_20_144_1": value  <=  3;
            "WIDTH_20_144_2": value  <=  3;
            "WIDTH_20_145_0": value  <=  4;
            "WIDTH_20_145_1": value  <=  2;
            "WIDTH_20_145_2": value  <=  2;
            "WIDTH_20_146_0": value  <=  2;
            "WIDTH_20_146_1": value  <=  1;
            "WIDTH_20_147_0": value  <=  3;
            "WIDTH_20_147_1": value  <=  1;
            "WIDTH_20_148_0": value  <=  3;
            "WIDTH_20_148_1": value  <=  1;
            "WIDTH_20_149_0": value  <=  4;
            "WIDTH_20_149_1": value  <=  2;
            "WIDTH_20_149_2": value  <=  2;
            "WIDTH_20_150_0": value  <=  4;
            "WIDTH_20_150_1": value  <=  2;
            "WIDTH_20_150_2": value  <=  2;
            "WIDTH_20_151_0": value  <=  2;
            "WIDTH_20_151_1": value  <=  1;
            "WIDTH_20_151_2": value  <=  1;
            "WIDTH_20_152_0": value  <=  2;
            "WIDTH_20_152_1": value  <=  1;
            "WIDTH_20_152_2": value  <=  1;
            "WIDTH_20_153_0": value  <=  6;
            "WIDTH_20_153_1": value  <=  6;
            "WIDTH_20_154_0": value  <=  12;
            "WIDTH_20_154_1": value  <=  4;
            "WIDTH_20_155_0": value  <=  3;
            "WIDTH_20_155_1": value  <=  1;
            "WIDTH_20_156_0": value  <=  3;
            "WIDTH_20_156_1": value  <=  1;
            "WIDTH_20_157_0": value  <=  6;
            "WIDTH_20_157_1": value  <=  6;
            "WIDTH_20_158_0": value  <=  3;
            "WIDTH_20_158_1": value  <=  1;
            "WIDTH_20_159_0": value  <=  6;
            "WIDTH_20_159_1": value  <=  3;
            "WIDTH_20_159_2": value  <=  3;
            "WIDTH_20_160_0": value  <=  6;
            "WIDTH_20_160_1": value  <=  2;
            "WIDTH_20_161_0": value  <=  2;
            "WIDTH_20_161_1": value  <=  1;
            "WIDTH_20_162_0": value  <=  8;
            "WIDTH_20_162_1": value  <=  4;
            "WIDTH_20_163_0": value  <=  8;
            "WIDTH_20_163_1": value  <=  8;
            "WIDTH_20_164_0": value  <=  4;
            "WIDTH_20_164_1": value  <=  4;
            "WIDTH_20_165_0": value  <=  4;
            "WIDTH_20_165_1": value  <=  4;
            "WIDTH_20_166_0": value  <=  17;
            "WIDTH_20_166_1": value  <=  17;
            "WIDTH_20_167_0": value  <=  4;
            "WIDTH_20_167_1": value  <=  4;
            "WIDTH_20_168_0": value  <=  6;
            "WIDTH_20_168_1": value  <=  6;
            "WIDTH_20_169_0": value  <=  5;
            "WIDTH_20_169_1": value  <=  5;
            "WIDTH_20_170_0": value  <=  2;
            "WIDTH_20_170_1": value  <=  1;
            "WIDTH_20_171_0": value  <=  2;
            "WIDTH_20_171_1": value  <=  1;
            "WIDTH_20_171_2": value  <=  1;
            "WIDTH_20_172_0": value  <=  11;
            "WIDTH_20_172_1": value  <=  11;
            "WIDTH_20_173_0": value  <=  6;
            "WIDTH_20_173_1": value  <=  3;
            "WIDTH_20_173_2": value  <=  3;
            "WIDTH_20_174_0": value  <=  4;
            "WIDTH_20_174_1": value  <=  4;
            "WIDTH_20_175_0": value  <=  3;
            "WIDTH_20_175_1": value  <=  1;
            "WIDTH_20_176_0": value  <=  3;
            "WIDTH_20_176_1": value  <=  3;
            "WIDTH_20_177_0": value  <=  2;
            "WIDTH_20_177_1": value  <=  2;
            "WIDTH_20_178_0": value  <=  16;
            "WIDTH_20_178_1": value  <=  16;
            "WIDTH_20_179_0": value  <=  2;
            "WIDTH_20_179_1": value  <=  1;
            "WIDTH_20_179_2": value  <=  1;
            "WIDTH_20_180_0": value  <=  2;
            "WIDTH_20_180_1": value  <=  1;
            "WIDTH_20_180_2": value  <=  1;
            "WIDTH_20_181_0": value  <=  3;
            "WIDTH_20_181_1": value  <=  3;
            "WIDTH_20_182_0": value  <=  3;
            "WIDTH_20_182_1": value  <=  3;
            "WIDTH_20_183_0": value  <=  10;
            "WIDTH_20_183_1": value  <=  5;
            "WIDTH_20_183_2": value  <=  5;
            "WIDTH_20_184_0": value  <=  14;
            "WIDTH_20_184_1": value  <=  14;
            "WIDTH_20_185_0": value  <=  1;
            "WIDTH_20_185_1": value  <=  1;
            "WIDTH_20_186_0": value  <=  2;
            "WIDTH_20_186_1": value  <=  1;
            "WIDTH_20_186_2": value  <=  1;
            "WIDTH_20_187_0": value  <=  2;
            "WIDTH_20_187_1": value  <=  2;
            "WIDTH_20_188_0": value  <=  20;
            "WIDTH_20_188_1": value  <=  10;
            "WIDTH_20_188_2": value  <=  10;
            "WIDTH_20_189_0": value  <=  1;
            "WIDTH_20_189_1": value  <=  1;
            "WIDTH_20_190_0": value  <=  3;
            "WIDTH_20_190_1": value  <=  1;
            "WIDTH_20_191_0": value  <=  3;
            "WIDTH_20_191_1": value  <=  1;
            "WIDTH_20_192_0": value  <=  2;
            "WIDTH_20_192_1": value  <=  1;
            "WIDTH_20_192_2": value  <=  1;
            "WIDTH_20_193_0": value  <=  3;
            "WIDTH_20_193_1": value  <=  1;
            "WIDTH_20_194_0": value  <=  1;
            "WIDTH_20_194_1": value  <=  1;
            "WIDTH_20_195_0": value  <=  5;
            "WIDTH_20_195_1": value  <=  5;
            "WIDTH_20_196_0": value  <=  6;
            "WIDTH_20_196_1": value  <=  3;
            "WIDTH_20_196_2": value  <=  3;
            "WIDTH_20_197_0": value  <=  3;
            "WIDTH_20_197_1": value  <=  1;
            "WIDTH_20_198_0": value  <=  12;
            "WIDTH_20_198_1": value  <=  4;
            "WIDTH_20_199_0": value  <=  5;
            "WIDTH_20_199_1": value  <=  5;
            "WIDTH_20_200_0": value  <=  14;
            "WIDTH_20_200_1": value  <=  7;
            "WIDTH_20_200_2": value  <=  7;
            "WIDTH_20_201_0": value  <=  14;
            "WIDTH_20_201_1": value  <=  7;
            "WIDTH_20_201_2": value  <=  7;
            "WIDTH_20_202_0": value  <=  4;
            "WIDTH_20_202_1": value  <=  4;
            "WIDTH_20_203_0": value  <=  6;
            "WIDTH_20_203_1": value  <=  2;
            "WIDTH_20_204_0": value  <=  1;
            "WIDTH_20_204_1": value  <=  1;
            "WIDTH_20_205_0": value  <=  6;
            "WIDTH_20_205_1": value  <=  2;
            "WIDTH_20_206_0": value  <=  3;
            "WIDTH_20_206_1": value  <=  1;
            "WIDTH_20_207_0": value  <=  9;
            "WIDTH_20_207_1": value  <=  9;
            "WIDTH_20_208_0": value  <=  20;
            "WIDTH_20_208_1": value  <=  10;
            "WIDTH_20_209_0": value  <=  4;
            "WIDTH_20_209_1": value  <=  2;
            "WIDTH_20_210_0": value  <=  2;
            "WIDTH_20_210_1": value  <=  2;
            "WIDTH_21_0_0": value  <=  10;
            "WIDTH_21_0_1": value  <=  10;
            "WIDTH_21_1_0": value  <=  4;
            "WIDTH_21_1_1": value  <=  2;
            "WIDTH_21_2_0": value  <=  2;
            "WIDTH_21_2_1": value  <=  1;
            "WIDTH_21_3_0": value  <=  12;
            "WIDTH_21_3_1": value  <=  4;
            "WIDTH_21_4_0": value  <=  9;
            "WIDTH_21_4_1": value  <=  3;
            "WIDTH_21_5_0": value  <=  1;
            "WIDTH_21_5_1": value  <=  1;
            "WIDTH_21_6_0": value  <=  6;
            "WIDTH_21_6_1": value  <=  3;
            "WIDTH_21_7_0": value  <=  1;
            "WIDTH_21_7_1": value  <=  1;
            "WIDTH_21_8_0": value  <=  6;
            "WIDTH_21_8_1": value  <=  6;
            "WIDTH_21_9_0": value  <=  2;
            "WIDTH_21_9_1": value  <=  1;
            "WIDTH_21_9_2": value  <=  1;
            "WIDTH_21_10_0": value  <=  1;
            "WIDTH_21_10_1": value  <=  1;
            "WIDTH_21_11_0": value  <=  5;
            "WIDTH_21_11_1": value  <=  5;
            "WIDTH_21_12_0": value  <=  4;
            "WIDTH_21_12_1": value  <=  2;
            "WIDTH_21_12_2": value  <=  2;
            "WIDTH_21_13_0": value  <=  16;
            "WIDTH_21_13_1": value  <=  8;
            "WIDTH_21_13_2": value  <=  8;
            "WIDTH_21_14_0": value  <=  1;
            "WIDTH_21_14_1": value  <=  1;
            "WIDTH_21_15_0": value  <=  15;
            "WIDTH_21_15_1": value  <=  5;
            "WIDTH_21_16_0": value  <=  15;
            "WIDTH_21_16_1": value  <=  5;
            "WIDTH_21_17_0": value  <=  3;
            "WIDTH_21_17_1": value  <=  3;
            "WIDTH_21_18_0": value  <=  8;
            "WIDTH_21_18_1": value  <=  4;
            "WIDTH_21_19_0": value  <=  2;
            "WIDTH_21_19_1": value  <=  2;
            "WIDTH_21_20_0": value  <=  16;
            "WIDTH_21_20_1": value  <=  16;
            "WIDTH_21_21_0": value  <=  7;
            "WIDTH_21_21_1": value  <=  7;
            "WIDTH_21_22_0": value  <=  10;
            "WIDTH_21_22_1": value  <=  10;
            "WIDTH_21_23_0": value  <=  3;
            "WIDTH_21_23_1": value  <=  1;
            "WIDTH_21_24_0": value  <=  1;
            "WIDTH_21_24_1": value  <=  1;
            "WIDTH_21_25_0": value  <=  14;
            "WIDTH_21_25_1": value  <=  14;
            "WIDTH_21_26_0": value  <=  3;
            "WIDTH_21_26_1": value  <=  1;
            "WIDTH_21_27_0": value  <=  5;
            "WIDTH_21_27_1": value  <=  5;
            "WIDTH_21_28_0": value  <=  5;
            "WIDTH_21_28_1": value  <=  5;
            "WIDTH_21_29_0": value  <=  2;
            "WIDTH_21_29_1": value  <=  2;
            "WIDTH_21_30_0": value  <=  2;
            "WIDTH_21_30_1": value  <=  2;
            "WIDTH_21_31_0": value  <=  2;
            "WIDTH_21_31_1": value  <=  2;
            "WIDTH_21_32_0": value  <=  2;
            "WIDTH_21_32_1": value  <=  2;
            "WIDTH_21_33_0": value  <=  10;
            "WIDTH_21_33_1": value  <=  5;
            "WIDTH_21_33_2": value  <=  5;
            "WIDTH_21_34_0": value  <=  1;
            "WIDTH_21_34_1": value  <=  1;
            "WIDTH_21_35_0": value  <=  2;
            "WIDTH_21_35_1": value  <=  1;
            "WIDTH_21_35_2": value  <=  1;
            "WIDTH_21_36_0": value  <=  2;
            "WIDTH_21_36_1": value  <=  2;
            "WIDTH_21_37_0": value  <=  6;
            "WIDTH_21_37_1": value  <=  6;
            "WIDTH_21_38_0": value  <=  2;
            "WIDTH_21_38_1": value  <=  2;
            "WIDTH_21_39_0": value  <=  4;
            "WIDTH_21_39_1": value  <=  4;
            "WIDTH_21_40_0": value  <=  4;
            "WIDTH_21_40_1": value  <=  4;
            "WIDTH_21_41_0": value  <=  2;
            "WIDTH_21_41_1": value  <=  1;
            "WIDTH_21_42_0": value  <=  8;
            "WIDTH_21_42_1": value  <=  4;
            "WIDTH_21_43_0": value  <=  4;
            "WIDTH_21_43_1": value  <=  4;
            "WIDTH_21_44_0": value  <=  10;
            "WIDTH_21_44_1": value  <=  10;
            "WIDTH_21_45_0": value  <=  1;
            "WIDTH_21_45_1": value  <=  1;
            "WIDTH_21_46_0": value  <=  4;
            "WIDTH_21_46_1": value  <=  4;
            "WIDTH_21_47_0": value  <=  8;
            "WIDTH_21_47_1": value  <=  4;
            "WIDTH_21_47_2": value  <=  4;
            "WIDTH_21_48_0": value  <=  4;
            "WIDTH_21_48_1": value  <=  2;
            "WIDTH_21_48_2": value  <=  2;
            "WIDTH_21_49_0": value  <=  3;
            "WIDTH_21_49_1": value  <=  1;
            "WIDTH_21_50_0": value  <=  2;
            "WIDTH_21_50_1": value  <=  1;
            "WIDTH_21_50_2": value  <=  1;
            "WIDTH_21_51_0": value  <=  6;
            "WIDTH_21_51_1": value  <=  2;
            "WIDTH_21_52_0": value  <=  2;
            "WIDTH_21_52_1": value  <=  2;
            "WIDTH_21_53_0": value  <=  1;
            "WIDTH_21_53_1": value  <=  1;
            "WIDTH_21_54_0": value  <=  6;
            "WIDTH_21_54_1": value  <=  3;
            "WIDTH_21_54_2": value  <=  3;
            "WIDTH_21_55_0": value  <=  3;
            "WIDTH_21_55_1": value  <=  1;
            "WIDTH_21_56_0": value  <=  2;
            "WIDTH_21_56_1": value  <=  2;
            "WIDTH_21_57_0": value  <=  3;
            "WIDTH_21_57_1": value  <=  1;
            "WIDTH_21_58_0": value  <=  3;
            "WIDTH_21_58_1": value  <=  3;
            "WIDTH_21_59_0": value  <=  2;
            "WIDTH_21_59_1": value  <=  1;
            "WIDTH_21_60_0": value  <=  18;
            "WIDTH_21_60_1": value  <=  6;
            "WIDTH_21_61_0": value  <=  4;
            "WIDTH_21_61_1": value  <=  2;
            "WIDTH_21_62_0": value  <=  4;
            "WIDTH_21_62_1": value  <=  2;
            "WIDTH_21_63_0": value  <=  2;
            "WIDTH_21_63_1": value  <=  1;
            "WIDTH_21_64_0": value  <=  2;
            "WIDTH_21_64_1": value  <=  1;
            "WIDTH_21_65_0": value  <=  2;
            "WIDTH_21_65_1": value  <=  1;
            "WIDTH_21_65_2": value  <=  1;
            "WIDTH_21_66_0": value  <=  2;
            "WIDTH_21_66_1": value  <=  1;
            "WIDTH_21_66_2": value  <=  1;
            "WIDTH_21_67_0": value  <=  3;
            "WIDTH_21_67_1": value  <=  1;
            "WIDTH_21_68_0": value  <=  3;
            "WIDTH_21_68_1": value  <=  3;
            "WIDTH_21_69_0": value  <=  4;
            "WIDTH_21_69_1": value  <=  4;
            "WIDTH_21_70_0": value  <=  3;
            "WIDTH_21_70_1": value  <=  1;
            "WIDTH_21_71_0": value  <=  3;
            "WIDTH_21_71_1": value  <=  1;
            "WIDTH_21_72_0": value  <=  3;
            "WIDTH_21_72_1": value  <=  1;
            "WIDTH_21_73_0": value  <=  3;
            "WIDTH_21_73_1": value  <=  1;
            "WIDTH_21_74_0": value  <=  3;
            "WIDTH_21_74_1": value  <=  1;
            "WIDTH_21_75_0": value  <=  12;
            "WIDTH_21_75_1": value  <=  6;
            "WIDTH_21_75_2": value  <=  6;
            "WIDTH_21_76_0": value  <=  2;
            "WIDTH_21_76_1": value  <=  2;
            "WIDTH_21_77_0": value  <=  3;
            "WIDTH_21_77_1": value  <=  3;
            "WIDTH_21_78_0": value  <=  4;
            "WIDTH_21_78_1": value  <=  2;
            "WIDTH_21_78_2": value  <=  2;
            "WIDTH_21_79_0": value  <=  3;
            "WIDTH_21_79_1": value  <=  1;
            "WIDTH_21_80_0": value  <=  1;
            "WIDTH_21_80_1": value  <=  1;
            "WIDTH_21_81_0": value  <=  3;
            "WIDTH_21_81_1": value  <=  1;
            "WIDTH_21_82_0": value  <=  3;
            "WIDTH_21_82_1": value  <=  1;
            "WIDTH_21_83_0": value  <=  15;
            "WIDTH_21_83_1": value  <=  15;
            "WIDTH_21_84_0": value  <=  2;
            "WIDTH_21_84_1": value  <=  1;
            "WIDTH_21_84_2": value  <=  1;
            "WIDTH_21_85_0": value  <=  2;
            "WIDTH_21_85_1": value  <=  2;
            "WIDTH_21_86_0": value  <=  3;
            "WIDTH_21_86_1": value  <=  1;
            "WIDTH_21_87_0": value  <=  3;
            "WIDTH_21_87_1": value  <=  3;
            "WIDTH_21_88_0": value  <=  3;
            "WIDTH_21_88_1": value  <=  3;
            "WIDTH_21_89_0": value  <=  6;
            "WIDTH_21_89_1": value  <=  3;
            "WIDTH_21_89_2": value  <=  3;
            "WIDTH_21_90_0": value  <=  12;
            "WIDTH_21_90_1": value  <=  4;
            "WIDTH_21_91_0": value  <=  2;
            "WIDTH_21_91_1": value  <=  2;
            "WIDTH_21_92_0": value  <=  1;
            "WIDTH_21_92_1": value  <=  1;
            "WIDTH_21_93_0": value  <=  6;
            "WIDTH_21_93_1": value  <=  3;
            "WIDTH_21_94_0": value  <=  3;
            "WIDTH_21_94_1": value  <=  1;
            "WIDTH_21_95_0": value  <=  2;
            "WIDTH_21_95_1": value  <=  1;
            "WIDTH_21_96_0": value  <=  2;
            "WIDTH_21_96_1": value  <=  1;
            "WIDTH_21_97_0": value  <=  2;
            "WIDTH_21_97_1": value  <=  1;
            "WIDTH_21_98_0": value  <=  10;
            "WIDTH_21_98_1": value  <=  5;
            "WIDTH_21_99_0": value  <=  3;
            "WIDTH_21_99_1": value  <=  1;
            "WIDTH_21_100_0": value  <=  9;
            "WIDTH_21_100_1": value  <=  3;
            "WIDTH_21_101_0": value  <=  2;
            "WIDTH_21_101_1": value  <=  2;
            "WIDTH_21_102_0": value  <=  16;
            "WIDTH_21_102_1": value  <=  8;
            "WIDTH_21_102_2": value  <=  8;
            "WIDTH_21_103_0": value  <=  2;
            "WIDTH_21_103_1": value  <=  1;
            "WIDTH_21_103_2": value  <=  1;
            "WIDTH_21_104_0": value  <=  2;
            "WIDTH_21_104_1": value  <=  2;
            "WIDTH_21_105_0": value  <=  3;
            "WIDTH_21_105_1": value  <=  1;
            "WIDTH_21_106_0": value  <=  8;
            "WIDTH_21_106_1": value  <=  8;
            "WIDTH_21_107_0": value  <=  2;
            "WIDTH_21_107_1": value  <=  2;
            "WIDTH_21_108_0": value  <=  2;
            "WIDTH_21_108_1": value  <=  2;
            "WIDTH_21_109_0": value  <=  3;
            "WIDTH_21_109_1": value  <=  3;
            "WIDTH_21_110_0": value  <=  2;
            "WIDTH_21_110_1": value  <=  2;
            "WIDTH_21_111_0": value  <=  3;
            "WIDTH_21_111_1": value  <=  3;
            "WIDTH_21_112_0": value  <=  3;
            "WIDTH_21_112_1": value  <=  3;
            "WIDTH_21_113_0": value  <=  2;
            "WIDTH_21_113_1": value  <=  1;
            "WIDTH_21_113_2": value  <=  1;
            "WIDTH_21_114_0": value  <=  3;
            "WIDTH_21_114_1": value  <=  1;
            "WIDTH_21_115_0": value  <=  6;
            "WIDTH_21_115_1": value  <=  2;
            "WIDTH_21_116_0": value  <=  6;
            "WIDTH_21_116_1": value  <=  2;
            "WIDTH_21_117_0": value  <=  1;
            "WIDTH_21_117_1": value  <=  1;
            "WIDTH_21_118_0": value  <=  10;
            "WIDTH_21_118_1": value  <=  10;
            "WIDTH_21_119_0": value  <=  1;
            "WIDTH_21_119_1": value  <=  1;
            "WIDTH_21_120_0": value  <=  2;
            "WIDTH_21_120_1": value  <=  1;
            "WIDTH_21_120_2": value  <=  1;
            "WIDTH_21_121_0": value  <=  2;
            "WIDTH_21_121_1": value  <=  1;
            "WIDTH_21_122_0": value  <=  1;
            "WIDTH_21_122_1": value  <=  1;
            "WIDTH_21_123_0": value  <=  3;
            "WIDTH_21_123_1": value  <=  1;
            "WIDTH_21_124_0": value  <=  2;
            "WIDTH_21_124_1": value  <=  1;
            "WIDTH_21_124_2": value  <=  1;
            "WIDTH_21_125_0": value  <=  3;
            "WIDTH_21_125_1": value  <=  1;
            "WIDTH_21_126_0": value  <=  3;
            "WIDTH_21_126_1": value  <=  1;
            "WIDTH_21_127_0": value  <=  8;
            "WIDTH_21_127_1": value  <=  4;
            "WIDTH_21_128_0": value  <=  8;
            "WIDTH_21_128_1": value  <=  4;
            "WIDTH_21_129_0": value  <=  2;
            "WIDTH_21_129_1": value  <=  1;
            "WIDTH_21_130_0": value  <=  2;
            "WIDTH_21_130_1": value  <=  1;
            "WIDTH_21_131_0": value  <=  2;
            "WIDTH_21_131_1": value  <=  2;
            "WIDTH_21_132_0": value  <=  3;
            "WIDTH_21_132_1": value  <=  3;
            "WIDTH_21_133_0": value  <=  1;
            "WIDTH_21_133_1": value  <=  1;
            "WIDTH_21_134_0": value  <=  18;
            "WIDTH_21_134_1": value  <=  9;
            "WIDTH_21_134_2": value  <=  9;
            "WIDTH_21_135_0": value  <=  1;
            "WIDTH_21_135_1": value  <=  1;
            "WIDTH_21_136_0": value  <=  2;
            "WIDTH_21_136_1": value  <=  2;
            "WIDTH_21_137_0": value  <=  3;
            "WIDTH_21_137_1": value  <=  1;
            "WIDTH_21_138_0": value  <=  18;
            "WIDTH_21_138_1": value  <=  18;
            "WIDTH_21_139_0": value  <=  14;
            "WIDTH_21_139_1": value  <=  14;
            "WIDTH_21_140_0": value  <=  3;
            "WIDTH_21_140_1": value  <=  1;
            "WIDTH_21_141_0": value  <=  3;
            "WIDTH_21_141_1": value  <=  1;
            "WIDTH_21_142_0": value  <=  1;
            "WIDTH_21_142_1": value  <=  1;
            "WIDTH_21_143_0": value  <=  6;
            "WIDTH_21_143_1": value  <=  6;
            "WIDTH_21_144_0": value  <=  7;
            "WIDTH_21_144_1": value  <=  7;
            "WIDTH_21_145_0": value  <=  6;
            "WIDTH_21_145_1": value  <=  6;
            "WIDTH_21_146_0": value  <=  6;
            "WIDTH_21_146_1": value  <=  2;
            "WIDTH_21_147_0": value  <=  6;
            "WIDTH_21_147_1": value  <=  3;
            "WIDTH_21_147_2": value  <=  3;
            "WIDTH_21_148_0": value  <=  18;
            "WIDTH_21_148_1": value  <=  18;
            "WIDTH_21_149_0": value  <=  17;
            "WIDTH_21_149_1": value  <=  17;
            "WIDTH_21_150_0": value  <=  7;
            "WIDTH_21_150_1": value  <=  7;
            "WIDTH_21_151_0": value  <=  1;
            "WIDTH_21_151_1": value  <=  1;
            "WIDTH_21_152_0": value  <=  3;
            "WIDTH_21_152_1": value  <=  3;
            "WIDTH_21_153_0": value  <=  6;
            "WIDTH_21_153_1": value  <=  6;
            "WIDTH_21_154_0": value  <=  6;
            "WIDTH_21_154_1": value  <=  6;
            "WIDTH_21_155_0": value  <=  4;
            "WIDTH_21_155_1": value  <=  4;
            "WIDTH_21_156_0": value  <=  4;
            "WIDTH_21_156_1": value  <=  4;
            "WIDTH_21_157_0": value  <=  2;
            "WIDTH_21_157_1": value  <=  2;
            "WIDTH_21_158_0": value  <=  4;
            "WIDTH_21_158_1": value  <=  2;
            "WIDTH_21_159_0": value  <=  8;
            "WIDTH_21_159_1": value  <=  4;
            "WIDTH_21_160_0": value  <=  4;
            "WIDTH_21_160_1": value  <=  2;
            "WIDTH_21_160_2": value  <=  2;
            "WIDTH_21_161_0": value  <=  2;
            "WIDTH_21_161_1": value  <=  2;
            "WIDTH_21_162_0": value  <=  1;
            "WIDTH_21_162_1": value  <=  1;
            "WIDTH_21_163_0": value  <=  2;
            "WIDTH_21_163_1": value  <=  2;
            "WIDTH_21_164_0": value  <=  4;
            "WIDTH_21_164_1": value  <=  4;
            "WIDTH_21_165_0": value  <=  8;
            "WIDTH_21_165_1": value  <=  8;
            "WIDTH_21_166_0": value  <=  6;
            "WIDTH_21_166_1": value  <=  3;
            "WIDTH_21_166_2": value  <=  3;
            "WIDTH_21_167_0": value  <=  3;
            "WIDTH_21_167_1": value  <=  1;
            "WIDTH_21_168_0": value  <=  2;
            "WIDTH_21_168_1": value  <=  2;
            "WIDTH_21_169_0": value  <=  6;
            "WIDTH_21_169_1": value  <=  6;
            "WIDTH_21_170_0": value  <=  19;
            "WIDTH_21_170_1": value  <=  19;
            "WIDTH_21_171_0": value  <=  8;
            "WIDTH_21_171_1": value  <=  8;
            "WIDTH_21_172_0": value  <=  3;
            "WIDTH_21_172_1": value  <=  1;
            "WIDTH_21_173_0": value  <=  4;
            "WIDTH_21_173_1": value  <=  2;
            "WIDTH_21_173_2": value  <=  2;
            "WIDTH_21_174_0": value  <=  6;
            "WIDTH_21_174_1": value  <=  6;
            "WIDTH_21_175_0": value  <=  4;
            "WIDTH_21_175_1": value  <=  4;
            "WIDTH_21_176_0": value  <=  3;
            "WIDTH_21_176_1": value  <=  1;
            "WIDTH_21_177_0": value  <=  3;
            "WIDTH_21_177_1": value  <=  1;
            "WIDTH_21_178_0": value  <=  3;
            "WIDTH_21_178_1": value  <=  1;
            "WIDTH_21_179_0": value  <=  6;
            "WIDTH_21_179_1": value  <=  2;
            "WIDTH_21_180_0": value  <=  4;
            "WIDTH_21_180_1": value  <=  2;
            "WIDTH_21_180_2": value  <=  2;
            "WIDTH_21_181_0": value  <=  4;
            "WIDTH_21_181_1": value  <=  2;
            "WIDTH_21_181_2": value  <=  2;
            "WIDTH_21_182_0": value  <=  1;
            "WIDTH_21_182_1": value  <=  1;
            "WIDTH_21_183_0": value  <=  2;
            "WIDTH_21_183_1": value  <=  1;
            "WIDTH_21_183_2": value  <=  1;
            "WIDTH_21_184_0": value  <=  2;
            "WIDTH_21_184_1": value  <=  1;
            "WIDTH_21_184_2": value  <=  1;
            "WIDTH_21_185_0": value  <=  14;
            "WIDTH_21_185_1": value  <=  14;
            "WIDTH_21_186_0": value  <=  3;
            "WIDTH_21_186_1": value  <=  3;
            "WIDTH_21_187_0": value  <=  2;
            "WIDTH_21_187_1": value  <=  2;
            "WIDTH_21_188_0": value  <=  6;
            "WIDTH_21_188_1": value  <=  6;
            "WIDTH_21_189_0": value  <=  3;
            "WIDTH_21_189_1": value  <=  3;
            "WIDTH_21_190_0": value  <=  3;
            "WIDTH_21_190_1": value  <=  3;
            "WIDTH_21_191_0": value  <=  2;
            "WIDTH_21_191_1": value  <=  2;
            "WIDTH_21_192_0": value  <=  18;
            "WIDTH_21_192_1": value  <=  6;
            "WIDTH_21_193_0": value  <=  6;
            "WIDTH_21_193_1": value  <=  6;
            "WIDTH_21_194_0": value  <=  18;
            "WIDTH_21_194_1": value  <=  6;
            "WIDTH_21_195_0": value  <=  2;
            "WIDTH_21_195_1": value  <=  1;
            "WIDTH_21_196_0": value  <=  2;
            "WIDTH_21_196_1": value  <=  1;
            "WIDTH_21_197_0": value  <=  2;
            "WIDTH_21_197_1": value  <=  2;
            "WIDTH_21_198_0": value  <=  3;
            "WIDTH_21_198_1": value  <=  1;
            "WIDTH_21_199_0": value  <=  3;
            "WIDTH_21_199_1": value  <=  1;
            "WIDTH_21_200_0": value  <=  3;
            "WIDTH_21_200_1": value  <=  1;
            "WIDTH_21_201_0": value  <=  3;
            "WIDTH_21_201_1": value  <=  1;
            "WIDTH_21_202_0": value  <=  3;
            "WIDTH_21_202_1": value  <=  1;
            "WIDTH_21_203_0": value  <=  6;
            "WIDTH_21_203_1": value  <=  6;
            "WIDTH_21_204_0": value  <=  2;
            "WIDTH_21_204_1": value  <=  2;
            "WIDTH_21_205_0": value  <=  1;
            "WIDTH_21_205_1": value  <=  1;
            "WIDTH_21_206_0": value  <=  8;
            "WIDTH_21_206_1": value  <=  4;
            "WIDTH_21_207_0": value  <=  20;
            "WIDTH_21_207_1": value  <=  10;
            "WIDTH_21_208_0": value  <=  1;
            "WIDTH_21_208_1": value  <=  1;
            "WIDTH_21_209_0": value  <=  4;
            "WIDTH_21_209_1": value  <=  4;
            "WIDTH_21_210_0": value  <=  14;
            "WIDTH_21_210_1": value  <=  14;
            "WIDTH_21_211_0": value  <=  18;
            "WIDTH_21_211_1": value  <=  18;
            "WIDTH_21_212_0": value  <=  10;
            "WIDTH_21_212_1": value  <=  5;
            "WIDTH_21_212_2": value  <=  5;

            default: value <= 0;

        endcase

    end

endmodule 
