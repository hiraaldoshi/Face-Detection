module Y_coord (

input string name,
output real value

);

always_comb
    begin

        case (name)

            Y_COORD_0_0_0: value  <=  7;
            Y_COORD_0_0_1: value  <=  9;
            Y_COORD_0_1_0: value  <=  2;
            Y_COORD_0_1_1: value  <=  2;
            Y_COORD_0_2_0: value  <=  7;
            Y_COORD_0_2_1: value  <=  10;
            Y_COORD_1_0_0: value  <=  6;
            Y_COORD_1_0_1: value  <=  9;
            Y_COORD_1_1_0: value  <=  5;
            Y_COORD_1_1_1: value  <=  5;
            Y_COORD_1_2_0: value  <=  0;
            Y_COORD_1_2_1: value  <=  3;
            Y_COORD_1_3_0: value  <=  9;
            Y_COORD_1_3_1: value  <=  13;
            Y_COORD_1_4_0: value  <=  6;
            Y_COORD_1_4_1: value  <=  10;
            Y_COORD_1_5_0: value  <=  1;
            Y_COORD_1_5_1: value  <=  1;
            Y_COORD_1_6_0: value  <=  8;
            Y_COORD_1_6_1: value  <=  12;
            Y_COORD_1_7_0: value  <=  1;
            Y_COORD_1_7_1: value  <=  1;
            Y_COORD_1_8_0: value  <=  8;
            Y_COORD_1_8_1: value  <=  9;
            Y_COORD_1_9_0: value  <=  6;
            Y_COORD_1_9_1: value  <=  7;
            Y_COORD_1_10_0: value  <=  17;
            Y_COORD_1_10_1: value  <=  18;
            Y_COORD_1_11_0: value  <=  2;
            Y_COORD_1_11_1: value  <=  2;
            Y_COORD_1_12_0: value  <=  0;
            Y_COORD_1_12_1: value  <=  0;
            Y_COORD_1_12_2: value  <=  6;
            Y_COORD_1_13_0: value  <=  11;
            Y_COORD_1_13_1: value  <=  11;
            Y_COORD_1_14_0: value  <=  7;
            Y_COORD_1_14_1: value  <=  8;
            Y_COORD_1_15_0: value  <=  11;
            Y_COORD_1_15_1: value  <=  12;
            Y_COORD_2_0_0: value  <=  3;
            Y_COORD_2_0_1: value  <=  6;
            Y_COORD_2_1_0: value  <=  4;
            Y_COORD_2_1_1: value  <=  11;
            Y_COORD_2_2_0: value  <=  5;
            Y_COORD_2_2_1: value  <=  9;
            Y_COORD_2_3_0: value  <=  5;
            Y_COORD_2_3_1: value  <=  5;
            Y_COORD_2_4_0: value  <=  6;
            Y_COORD_2_4_1: value  <=  10;
            Y_COORD_2_5_0: value  <=  0;
            Y_COORD_2_5_1: value  <=  3;
            Y_COORD_2_6_0: value  <=  12;
            Y_COORD_2_6_1: value  <=  16;
            Y_COORD_2_7_0: value  <=  7;
            Y_COORD_2_7_1: value  <=  9;
            Y_COORD_2_8_0: value  <=  0;
            Y_COORD_2_8_1: value  <=  0;
            Y_COORD_2_9_0: value  <=  0;
            Y_COORD_2_9_1: value  <=  0;
            Y_COORD_2_10_0: value  <=  1;
            Y_COORD_2_10_1: value  <=  1;
            Y_COORD_2_11_0: value  <=  1;
            Y_COORD_2_11_1: value  <=  1;
            Y_COORD_2_12_0: value  <=  5;
            Y_COORD_2_12_1: value  <=  5;
            Y_COORD_2_12_2: value  <=  9;
            Y_COORD_2_13_0: value  <=  15;
            Y_COORD_2_13_1: value  <=  15;
            Y_COORD_2_13_2: value  <=  17;
            Y_COORD_2_14_0: value  <=  1;
            Y_COORD_2_14_1: value  <=  1;
            Y_COORD_2_14_2: value  <=  5;
            Y_COORD_2_15_0: value  <=  6;
            Y_COORD_2_15_1: value  <=  6;
            Y_COORD_2_15_2: value  <=  11;
            Y_COORD_2_16_0: value  <=  1;
            Y_COORD_2_16_1: value  <=  1;
            Y_COORD_2_17_0: value  <=  18;
            Y_COORD_2_17_1: value  <=  19;
            Y_COORD_2_18_0: value  <=  13;
            Y_COORD_2_18_1: value  <=  14;
            Y_COORD_2_19_0: value  <=  14;
            Y_COORD_2_19_1: value  <=  15;
            Y_COORD_2_20_0: value  <=  12;
            Y_COORD_2_20_1: value  <=  14;
            Y_COORD_3_0_0: value  <=  7;
            Y_COORD_3_0_1: value  <=  9;
            Y_COORD_3_1_0: value  <=  3;
            Y_COORD_3_1_1: value  <=  11;
            Y_COORD_3_2_0: value  <=  6;
            Y_COORD_3_2_1: value  <=  10;
            Y_COORD_3_3_0: value  <=  3;
            Y_COORD_3_3_1: value  <=  3;
            Y_COORD_3_4_0: value  <=  8;
            Y_COORD_3_4_1: value  <=  12;
            Y_COORD_3_5_0: value  <=  3;
            Y_COORD_3_5_1: value  <=  3;
            Y_COORD_3_5_2: value  <=  6;
            Y_COORD_3_6_0: value  <=  1;
            Y_COORD_3_6_1: value  <=  1;
            Y_COORD_3_7_0: value  <=  0;
            Y_COORD_3_7_1: value  <=  0;
            Y_COORD_3_8_0: value  <=  1;
            Y_COORD_3_8_1: value  <=  1;
            Y_COORD_3_9_0: value  <=  15;
            Y_COORD_3_9_1: value  <=  15;
            Y_COORD_3_9_2: value  <=  17;
            Y_COORD_3_10_0: value  <=  3;
            Y_COORD_3_10_1: value  <=  3;
            Y_COORD_3_11_0: value  <=  4;
            Y_COORD_3_11_1: value  <=  9;
            Y_COORD_3_12_0: value  <=  5;
            Y_COORD_3_12_1: value  <=  7;
            Y_COORD_3_13_0: value  <=  4;
            Y_COORD_3_13_1: value  <=  4;
            Y_COORD_3_13_2: value  <=  9;
            Y_COORD_3_14_0: value  <=  4;
            Y_COORD_3_14_1: value  <=  4;
            Y_COORD_3_15_0: value  <=  11;
            Y_COORD_3_15_1: value  <=  12;
            Y_COORD_3_16_0: value  <=  11;
            Y_COORD_3_16_1: value  <=  12;
            Y_COORD_3_17_0: value  <=  11;
            Y_COORD_3_17_1: value  <=  12;
            Y_COORD_3_18_0: value  <=  15;
            Y_COORD_3_18_1: value  <=  15;
            Y_COORD_3_18_2: value  <=  17;
            Y_COORD_3_19_0: value  <=  7;
            Y_COORD_3_19_1: value  <=  8;
            Y_COORD_3_20_0: value  <=  11;
            Y_COORD_3_20_1: value  <=  12;
            Y_COORD_3_21_0: value  <=  0;
            Y_COORD_3_21_1: value  <=  1;
            Y_COORD_3_22_0: value  <=  14;
            Y_COORD_3_22_1: value  <=  15;
            Y_COORD_3_23_0: value  <=  15;
            Y_COORD_3_23_1: value  <=  16;
            Y_COORD_3_24_0: value  <=  5;
            Y_COORD_3_24_1: value  <=  7;
            Y_COORD_3_25_0: value  <=  12;
            Y_COORD_3_25_1: value  <=  12;
            Y_COORD_3_26_0: value  <=  3;
            Y_COORD_3_26_1: value  <=  6;
            Y_COORD_3_27_0: value  <=  17;
            Y_COORD_3_27_1: value  <=  17;
            Y_COORD_3_28_0: value  <=  9;
            Y_COORD_3_28_1: value  <=  10;
            Y_COORD_3_29_0: value  <=  6;
            Y_COORD_3_29_1: value  <=  6;
            Y_COORD_3_30_0: value  <=  17;
            Y_COORD_3_30_1: value  <=  17;
            Y_COORD_3_31_0: value  <=  17;
            Y_COORD_3_31_1: value  <=  17;
            Y_COORD_3_32_0: value  <=  12;
            Y_COORD_3_32_1: value  <=  13;
            Y_COORD_3_33_0: value  <=  3;
            Y_COORD_3_33_1: value  <=  3;
            Y_COORD_3_34_0: value  <=  11;
            Y_COORD_3_34_1: value  <=  13;
            Y_COORD_3_35_0: value  <=  10;
            Y_COORD_3_35_1: value  <=  10;
            Y_COORD_3_35_2: value  <=  12;
            Y_COORD_3_36_0: value  <=  10;
            Y_COORD_3_36_1: value  <=  11;
            Y_COORD_3_37_0: value  <=  1;
            Y_COORD_3_37_1: value  <=  1;
            Y_COORD_3_38_0: value  <=  7;
            Y_COORD_3_38_1: value  <=  7;
            Y_COORD_4_0_0: value  <=  0;
            Y_COORD_4_0_1: value  <=  3;
            Y_COORD_4_1_0: value  <=  10;
            Y_COORD_4_1_1: value  <=  13;
            Y_COORD_4_2_0: value  <=  5;
            Y_COORD_4_2_1: value  <=  9;
            Y_COORD_4_3_0: value  <=  0;
            Y_COORD_4_3_1: value  <=  0;
            Y_COORD_4_4_0: value  <=  3;
            Y_COORD_4_4_1: value  <=  3;
            Y_COORD_4_5_0: value  <=  3;
            Y_COORD_4_5_1: value  <=  3;
            Y_COORD_4_6_0: value  <=  10;
            Y_COORD_4_6_1: value  <=  13;
            Y_COORD_4_7_0: value  <=  3;
            Y_COORD_4_7_1: value  <=  3;
            Y_COORD_4_8_0: value  <=  4;
            Y_COORD_4_8_1: value  <=  6;
            Y_COORD_4_9_0: value  <=  12;
            Y_COORD_4_9_1: value  <=  14;
            Y_COORD_4_10_0: value  <=  3;
            Y_COORD_4_10_1: value  <=  3;
            Y_COORD_4_11_0: value  <=  3;
            Y_COORD_4_11_1: value  <=  3;
            Y_COORD_4_12_0: value  <=  1;
            Y_COORD_4_12_1: value  <=  1;
            Y_COORD_4_13_0: value  <=  0;
            Y_COORD_4_13_1: value  <=  0;
            Y_COORD_4_13_2: value  <=  2;
            Y_COORD_4_14_0: value  <=  5;
            Y_COORD_4_14_1: value  <=  12;
            Y_COORD_4_15_0: value  <=  0;
            Y_COORD_4_15_1: value  <=  2;
            Y_COORD_4_16_0: value  <=  5;
            Y_COORD_4_16_1: value  <=  5;
            Y_COORD_4_17_0: value  <=  18;
            Y_COORD_4_17_1: value  <=  18;
            Y_COORD_4_18_0: value  <=  18;
            Y_COORD_4_18_1: value  <=  18;
            Y_COORD_4_19_0: value  <=  5;
            Y_COORD_4_19_1: value  <=  7;
            Y_COORD_4_20_0: value  <=  12;
            Y_COORD_4_20_1: value  <=  14;
            Y_COORD_4_21_0: value  <=  8;
            Y_COORD_4_21_1: value  <=  12;
            Y_COORD_4_22_0: value  <=  18;
            Y_COORD_4_22_1: value  <=  18;
            Y_COORD_4_23_0: value  <=  0;
            Y_COORD_4_23_1: value  <=  0;
            Y_COORD_4_24_0: value  <=  11;
            Y_COORD_4_24_1: value  <=  12;
            Y_COORD_4_25_0: value  <=  0;
            Y_COORD_4_25_1: value  <=  0;
            Y_COORD_4_26_0: value  <=  1;
            Y_COORD_4_26_1: value  <=  1;
            Y_COORD_4_27_0: value  <=  0;
            Y_COORD_4_27_1: value  <=  0;
            Y_COORD_4_27_2: value  <=  2;
            Y_COORD_4_28_0: value  <=  12;
            Y_COORD_4_28_1: value  <=  13;
            Y_COORD_4_29_0: value  <=  14;
            Y_COORD_4_29_1: value  <=  15;
            Y_COORD_4_30_0: value  <=  4;
            Y_COORD_4_30_1: value  <=  4;
            Y_COORD_4_30_2: value  <=  10;
            Y_COORD_4_31_0: value  <=  6;
            Y_COORD_4_31_1: value  <=  10;
            Y_COORD_4_32_0: value  <=  2;
            Y_COORD_4_32_1: value  <=  2;
            Y_COORD_4_32_2: value  <=  9;
            Y_COORD_5_0_0: value  <=  7;
            Y_COORD_5_0_1: value  <=  7;
            Y_COORD_5_1_0: value  <=  4;
            Y_COORD_5_1_1: value  <=  6;
            Y_COORD_5_2_0: value  <=  5;
            Y_COORD_5_2_1: value  <=  9;
            Y_COORD_5_3_0: value  <=  10;
            Y_COORD_5_3_1: value  <=  12;
            Y_COORD_5_4_0: value  <=  0;
            Y_COORD_5_4_1: value  <=  1;
            Y_COORD_5_5_0: value  <=  5;
            Y_COORD_5_5_1: value  <=  5;
            Y_COORD_5_6_0: value  <=  2;
            Y_COORD_5_6_1: value  <=  2;
            Y_COORD_5_6_2: value  <=  7;
            Y_COORD_5_7_0: value  <=  5;
            Y_COORD_5_7_1: value  <=  10;
            Y_COORD_5_8_0: value  <=  14;
            Y_COORD_5_8_1: value  <=  14;
            Y_COORD_5_8_2: value  <=  17;
            Y_COORD_5_9_0: value  <=  2;
            Y_COORD_5_9_1: value  <=  3;
            Y_COORD_5_10_0: value  <=  10;
            Y_COORD_5_10_1: value  <=  13;
            Y_COORD_5_11_0: value  <=  4;
            Y_COORD_5_11_1: value  <=  4;
            Y_COORD_5_12_0: value  <=  9;
            Y_COORD_5_12_1: value  <=  9;
            Y_COORD_5_12_2: value  <=  12;
            Y_COORD_5_13_0: value  <=  7;
            Y_COORD_5_13_1: value  <=  9;
            Y_COORD_5_14_0: value  <=  9;
            Y_COORD_5_14_1: value  <=  9;
            Y_COORD_5_14_2: value  <=  13;
            Y_COORD_5_15_0: value  <=  1;
            Y_COORD_5_15_1: value  <=  2;
            Y_COORD_5_16_0: value  <=  4;
            Y_COORD_5_16_1: value  <=  4;
            Y_COORD_5_17_0: value  <=  10;
            Y_COORD_5_17_1: value  <=  14;
            Y_COORD_5_18_0: value  <=  0;
            Y_COORD_5_18_1: value  <=  1;
            Y_COORD_5_19_0: value  <=  5;
            Y_COORD_5_19_1: value  <=  5;
            Y_COORD_5_19_2: value  <=  9;
            Y_COORD_5_20_0: value  <=  6;
            Y_COORD_5_20_1: value  <=  9;
            Y_COORD_5_21_0: value  <=  1;
            Y_COORD_5_21_1: value  <=  2;
            Y_COORD_5_22_0: value  <=  6;
            Y_COORD_5_22_1: value  <=  6;
            Y_COORD_5_23_0: value  <=  1;
            Y_COORD_5_23_1: value  <=  2;
            Y_COORD_5_24_0: value  <=  13;
            Y_COORD_5_24_1: value  <=  14;
            Y_COORD_5_25_0: value  <=  4;
            Y_COORD_5_25_1: value  <=  4;
            Y_COORD_5_25_2: value  <=  10;
            Y_COORD_5_26_0: value  <=  2;
            Y_COORD_5_26_1: value  <=  2;
            Y_COORD_5_27_0: value  <=  1;
            Y_COORD_5_27_1: value  <=  6;
            Y_COORD_5_28_0: value  <=  4;
            Y_COORD_5_28_1: value  <=  4;
            Y_COORD_5_29_0: value  <=  13;
            Y_COORD_5_29_1: value  <=  14;
            Y_COORD_5_30_0: value  <=  14;
            Y_COORD_5_30_1: value  <=  15;
            Y_COORD_5_31_0: value  <=  13;
            Y_COORD_5_31_1: value  <=  14;
            Y_COORD_5_32_0: value  <=  14;
            Y_COORD_5_32_1: value  <=  15;
            Y_COORD_5_33_0: value  <=  13;
            Y_COORD_5_33_1: value  <=  14;
            Y_COORD_5_34_0: value  <=  13;
            Y_COORD_5_34_1: value  <=  14;
            Y_COORD_5_35_0: value  <=  7;
            Y_COORD_5_35_1: value  <=  7;
            Y_COORD_5_35_2: value  <=  13;
            Y_COORD_5_36_0: value  <=  7;
            Y_COORD_5_36_1: value  <=  7;
            Y_COORD_5_37_0: value  <=  9;
            Y_COORD_5_37_1: value  <=  10;
            Y_COORD_5_38_0: value  <=  6;
            Y_COORD_5_38_1: value  <=  6;
            Y_COORD_5_39_0: value  <=  6;
            Y_COORD_5_39_1: value  <=  10;
            Y_COORD_5_40_0: value  <=  7;
            Y_COORD_5_40_1: value  <=  7;
            Y_COORD_5_41_0: value  <=  3;
            Y_COORD_5_41_1: value  <=  3;
            Y_COORD_5_42_0: value  <=  4;
            Y_COORD_5_42_1: value  <=  4;
            Y_COORD_5_43_0: value  <=  6;
            Y_COORD_5_43_1: value  <=  7;
            Y_COORD_6_0_0: value  <=  3;
            Y_COORD_6_0_1: value  <=  6;
            Y_COORD_6_1_0: value  <=  7;
            Y_COORD_6_1_1: value  <=  7;
            Y_COORD_6_2_0: value  <=  8;
            Y_COORD_6_2_1: value  <=  12;
            Y_COORD_6_3_0: value  <=  6;
            Y_COORD_6_3_1: value  <=  9;
            Y_COORD_6_4_0: value  <=  5;
            Y_COORD_6_4_1: value  <=  10;
            Y_COORD_6_5_0: value  <=  0;
            Y_COORD_6_5_1: value  <=  3;
            Y_COORD_6_6_0: value  <=  6;
            Y_COORD_6_6_1: value  <=  13;
            Y_COORD_6_7_0: value  <=  7;
            Y_COORD_6_7_1: value  <=  9;
            Y_COORD_6_8_0: value  <=  8;
            Y_COORD_6_8_1: value  <=  8;
            Y_COORD_6_9_0: value  <=  2;
            Y_COORD_6_9_1: value  <=  7;
            Y_COORD_6_10_0: value  <=  7;
            Y_COORD_6_10_1: value  <=  9;
            Y_COORD_6_11_0: value  <=  3;
            Y_COORD_6_11_1: value  <=  3;
            Y_COORD_6_12_0: value  <=  7;
            Y_COORD_6_12_1: value  <=  7;
            Y_COORD_6_12_2: value  <=  12;
            Y_COORD_6_13_0: value  <=  4;
            Y_COORD_6_13_1: value  <=  4;
            Y_COORD_6_13_2: value  <=  10;
            Y_COORD_6_14_0: value  <=  4;
            Y_COORD_6_14_1: value  <=  4;
            Y_COORD_6_15_0: value  <=  3;
            Y_COORD_6_15_1: value  <=  3;
            Y_COORD_6_16_0: value  <=  3;
            Y_COORD_6_16_1: value  <=  3;
            Y_COORD_6_17_0: value  <=  14;
            Y_COORD_6_17_1: value  <=  15;
            Y_COORD_6_18_0: value  <=  12;
            Y_COORD_6_18_1: value  <=  12;
            Y_COORD_6_19_0: value  <=  14;
            Y_COORD_6_19_1: value  <=  15;
            Y_COORD_6_20_0: value  <=  11;
            Y_COORD_6_20_1: value  <=  14;
            Y_COORD_6_21_0: value  <=  11;
            Y_COORD_6_21_1: value  <=  14;
            Y_COORD_6_22_0: value  <=  15;
            Y_COORD_6_22_1: value  <=  16;
            Y_COORD_6_23_0: value  <=  0;
            Y_COORD_6_23_1: value  <=  0;
            Y_COORD_6_24_0: value  <=  5;
            Y_COORD_6_24_1: value  <=  5;
            Y_COORD_6_25_0: value  <=  0;
            Y_COORD_6_25_1: value  <=  3;
            Y_COORD_6_26_0: value  <=  2;
            Y_COORD_6_26_1: value  <=  2;
            Y_COORD_6_26_2: value  <=  6;
            Y_COORD_6_27_0: value  <=  12;
            Y_COORD_6_27_1: value  <=  14;
            Y_COORD_6_28_0: value  <=  12;
            Y_COORD_6_28_1: value  <=  14;
            Y_COORD_6_29_0: value  <=  11;
            Y_COORD_6_29_1: value  <=  13;
            Y_COORD_6_30_0: value  <=  4;
            Y_COORD_6_30_1: value  <=  5;
            Y_COORD_6_31_0: value  <=  5;
            Y_COORD_6_31_1: value  <=  9;
            Y_COORD_6_32_0: value  <=  8;
            Y_COORD_6_32_1: value  <=  8;
            Y_COORD_6_33_0: value  <=  1;
            Y_COORD_6_33_1: value  <=  1;
            Y_COORD_6_34_0: value  <=  5;
            Y_COORD_6_34_1: value  <=  6;
            Y_COORD_6_35_0: value  <=  9;
            Y_COORD_6_35_1: value  <=  9;
            Y_COORD_6_35_2: value  <=  12;
            Y_COORD_6_36_0: value  <=  6;
            Y_COORD_6_36_1: value  <=  6;
            Y_COORD_6_37_0: value  <=  0;
            Y_COORD_6_37_1: value  <=  1;
            Y_COORD_6_38_0: value  <=  2;
            Y_COORD_6_38_1: value  <=  3;
            Y_COORD_6_39_0: value  <=  6;
            Y_COORD_6_39_1: value  <=  7;
            Y_COORD_6_40_0: value  <=  0;
            Y_COORD_6_40_1: value  <=  0;
            Y_COORD_6_41_0: value  <=  7;
            Y_COORD_6_41_1: value  <=  7;
            Y_COORD_6_42_0: value  <=  7;
            Y_COORD_6_42_1: value  <=  7;
            Y_COORD_6_43_0: value  <=  7;
            Y_COORD_6_43_1: value  <=  7;
            Y_COORD_6_43_2: value  <=  9;
            Y_COORD_6_44_0: value  <=  5;
            Y_COORD_6_44_1: value  <=  7;
            Y_COORD_6_45_0: value  <=  11;
            Y_COORD_6_45_1: value  <=  13;
            Y_COORD_6_46_0: value  <=  11;
            Y_COORD_6_46_1: value  <=  13;
            Y_COORD_6_47_0: value  <=  9;
            Y_COORD_6_47_1: value  <=  9;
            Y_COORD_6_47_2: value  <=  13;
            Y_COORD_6_48_0: value  <=  12;
            Y_COORD_6_48_1: value  <=  13;
            Y_COORD_6_49_0: value  <=  15;
            Y_COORD_6_49_1: value  <=  17;
            Y_COORD_7_0_0: value  <=  7;
            Y_COORD_7_0_1: value  <=  7;
            Y_COORD_7_1_0: value  <=  3;
            Y_COORD_7_1_1: value  <=  3;
            Y_COORD_7_1_2: value  <=  6;
            Y_COORD_7_2_0: value  <=  4;
            Y_COORD_7_2_1: value  <=  6;
            Y_COORD_7_3_0: value  <=  3;
            Y_COORD_7_3_1: value  <=  3;
            Y_COORD_7_3_2: value  <=  10;
            Y_COORD_7_4_0: value  <=  4;
            Y_COORD_7_4_1: value  <=  9;
            Y_COORD_7_5_0: value  <=  2;
            Y_COORD_7_5_1: value  <=  2;
            Y_COORD_7_5_2: value  <=  6;
            Y_COORD_7_6_0: value  <=  2;
            Y_COORD_7_6_1: value  <=  2;
            Y_COORD_7_6_2: value  <=  6;
            Y_COORD_7_7_0: value  <=  13;
            Y_COORD_7_7_1: value  <=  13;
            Y_COORD_7_8_0: value  <=  3;
            Y_COORD_7_8_1: value  <=  3;
            Y_COORD_7_8_2: value  <=  10;
            Y_COORD_7_9_0: value  <=  1;
            Y_COORD_7_9_1: value  <=  3;
            Y_COORD_7_10_0: value  <=  11;
            Y_COORD_7_10_1: value  <=  12;
            Y_COORD_7_11_0: value  <=  1;
            Y_COORD_7_11_1: value  <=  3;
            Y_COORD_7_12_0: value  <=  1;
            Y_COORD_7_12_1: value  <=  3;
            Y_COORD_7_13_0: value  <=  5;
            Y_COORD_7_13_1: value  <=  7;
            Y_COORD_7_14_0: value  <=  2;
            Y_COORD_7_14_1: value  <=  2;
            Y_COORD_7_15_0: value  <=  3;
            Y_COORD_7_15_1: value  <=  10;
            Y_COORD_7_16_0: value  <=  7;
            Y_COORD_7_16_1: value  <=  12;
            Y_COORD_7_17_0: value  <=  15;
            Y_COORD_7_17_1: value  <=  16;
            Y_COORD_7_18_0: value  <=  11;
            Y_COORD_7_18_1: value  <=  11;
            Y_COORD_7_18_2: value  <=  13;
            Y_COORD_7_19_0: value  <=  7;
            Y_COORD_7_19_1: value  <=  7;
            Y_COORD_7_19_2: value  <=  9;
            Y_COORD_7_20_0: value  <=  10;
            Y_COORD_7_20_1: value  <=  13;
            Y_COORD_7_21_0: value  <=  6;
            Y_COORD_7_21_1: value  <=  9;
            Y_COORD_7_22_0: value  <=  10;
            Y_COORD_7_22_1: value  <=  10;
            Y_COORD_7_23_0: value  <=  8;
            Y_COORD_7_23_1: value  <=  8;
            Y_COORD_7_24_0: value  <=  6;
            Y_COORD_7_24_1: value  <=  8;
            Y_COORD_7_25_0: value  <=  1;
            Y_COORD_7_25_1: value  <=  3;
            Y_COORD_7_26_0: value  <=  7;
            Y_COORD_7_26_1: value  <=  7;
            Y_COORD_7_27_0: value  <=  7;
            Y_COORD_7_27_1: value  <=  7;
            Y_COORD_7_28_0: value  <=  7;
            Y_COORD_7_28_1: value  <=  7;
            Y_COORD_7_29_0: value  <=  9;
            Y_COORD_7_29_1: value  <=  10;
            Y_COORD_7_30_0: value  <=  8;
            Y_COORD_7_30_1: value  <=  9;
            Y_COORD_7_31_0: value  <=  5;
            Y_COORD_7_31_1: value  <=  5;
            Y_COORD_7_32_0: value  <=  13;
            Y_COORD_7_32_1: value  <=  14;
            Y_COORD_7_33_0: value  <=  7;
            Y_COORD_7_33_1: value  <=  7;
            Y_COORD_7_33_2: value  <=  10;
            Y_COORD_7_34_0: value  <=  14;
            Y_COORD_7_34_1: value  <=  15;
            Y_COORD_7_35_0: value  <=  7;
            Y_COORD_7_35_1: value  <=  8;
            Y_COORD_7_36_0: value  <=  4;
            Y_COORD_7_36_1: value  <=  4;
            Y_COORD_7_37_0: value  <=  0;
            Y_COORD_7_37_1: value  <=  0;
            Y_COORD_7_38_0: value  <=  3;
            Y_COORD_7_38_1: value  <=  3;
            Y_COORD_7_39_0: value  <=  3;
            Y_COORD_7_39_1: value  <=  3;
            Y_COORD_7_40_0: value  <=  13;
            Y_COORD_7_40_1: value  <=  16;
            Y_COORD_7_41_0: value  <=  3;
            Y_COORD_7_41_1: value  <=  3;
            Y_COORD_7_42_0: value  <=  7;
            Y_COORD_7_42_1: value  <=  7;
            Y_COORD_7_42_2: value  <=  9;
            Y_COORD_7_43_0: value  <=  3;
            Y_COORD_7_43_1: value  <=  3;
            Y_COORD_7_44_0: value  <=  3;
            Y_COORD_7_44_1: value  <=  3;
            Y_COORD_7_45_0: value  <=  1;
            Y_COORD_7_45_1: value  <=  1;
            Y_COORD_7_46_0: value  <=  0;
            Y_COORD_7_46_1: value  <=  0;
            Y_COORD_7_47_0: value  <=  16;
            Y_COORD_7_47_1: value  <=  16;
            Y_COORD_7_47_2: value  <=  18;
            Y_COORD_7_48_0: value  <=  6;
            Y_COORD_7_48_1: value  <=  6;
            Y_COORD_7_49_0: value  <=  5;
            Y_COORD_7_49_1: value  <=  5;
            Y_COORD_7_50_0: value  <=  7;
            Y_COORD_7_50_1: value  <=  7;
            Y_COORD_8_0_0: value  <=  4;
            Y_COORD_8_0_1: value  <=  6;
            Y_COORD_8_1_0: value  <=  5;
            Y_COORD_8_1_1: value  <=  11;
            Y_COORD_8_2_0: value  <=  6;
            Y_COORD_8_2_1: value  <=  10;
            Y_COORD_8_3_0: value  <=  2;
            Y_COORD_8_3_1: value  <=  2;
            Y_COORD_8_4_0: value  <=  8;
            Y_COORD_8_4_1: value  <=  9;
            Y_COORD_8_5_0: value  <=  12;
            Y_COORD_8_5_1: value  <=  16;
            Y_COORD_8_6_0: value  <=  2;
            Y_COORD_8_6_1: value  <=  2;
            Y_COORD_8_7_0: value  <=  11;
            Y_COORD_8_7_1: value  <=  13;
            Y_COORD_8_8_0: value  <=  11;
            Y_COORD_8_8_1: value  <=  11;
            Y_COORD_8_9_0: value  <=  3;
            Y_COORD_8_9_1: value  <=  3;
            Y_COORD_8_10_0: value  <=  13;
            Y_COORD_8_10_1: value  <=  14;
            Y_COORD_8_11_0: value  <=  11;
            Y_COORD_8_11_1: value  <=  14;
            Y_COORD_8_12_0: value  <=  11;
            Y_COORD_8_12_1: value  <=  14;
            Y_COORD_8_13_0: value  <=  14;
            Y_COORD_8_13_1: value  <=  16;
            Y_COORD_8_14_0: value  <=  14;
            Y_COORD_8_14_1: value  <=  15;
            Y_COORD_8_15_0: value  <=  0;
            Y_COORD_8_15_1: value  <=  0;
            Y_COORD_8_16_0: value  <=  1;
            Y_COORD_8_16_1: value  <=  1;
            Y_COORD_8_17_0: value  <=  3;
            Y_COORD_8_17_1: value  <=  3;
            Y_COORD_8_18_0: value  <=  8;
            Y_COORD_8_18_1: value  <=  10;
            Y_COORD_8_19_0: value  <=  12;
            Y_COORD_8_19_1: value  <=  13;
            Y_COORD_8_20_0: value  <=  18;
            Y_COORD_8_20_1: value  <=  19;
            Y_COORD_8_21_0: value  <=  1;
            Y_COORD_8_21_1: value  <=  3;
            Y_COORD_8_22_0: value  <=  0;
            Y_COORD_8_22_1: value  <=  0;
            Y_COORD_8_23_0: value  <=  8;
            Y_COORD_8_23_1: value  <=  8;
            Y_COORD_8_23_2: value  <=  9;
            Y_COORD_8_24_0: value  <=  10;
            Y_COORD_8_24_1: value  <=  13;
            Y_COORD_8_25_0: value  <=  13;
            Y_COORD_8_25_1: value  <=  13;
            Y_COORD_8_25_2: value  <=  15;
            Y_COORD_8_26_0: value  <=  7;
            Y_COORD_8_26_1: value  <=  7;
            Y_COORD_8_27_0: value  <=  0;
            Y_COORD_8_27_1: value  <=  1;
            Y_COORD_8_28_0: value  <=  8;
            Y_COORD_8_28_1: value  <=  8;
            Y_COORD_8_28_2: value  <=  9;
            Y_COORD_8_29_0: value  <=  2;
            Y_COORD_8_29_1: value  <=  2;
            Y_COORD_8_29_2: value  <=  3;
            Y_COORD_8_30_0: value  <=  14;
            Y_COORD_8_30_1: value  <=  15;
            Y_COORD_8_31_0: value  <=  13;
            Y_COORD_8_31_1: value  <=  13;
            Y_COORD_8_31_2: value  <=  16;
            Y_COORD_8_32_0: value  <=  12;
            Y_COORD_8_32_1: value  <=  13;
            Y_COORD_8_33_0: value  <=  11;
            Y_COORD_8_33_1: value  <=  13;
            Y_COORD_8_34_0: value  <=  11;
            Y_COORD_8_34_1: value  <=  13;
            Y_COORD_8_35_0: value  <=  4;
            Y_COORD_8_35_1: value  <=  4;
            Y_COORD_8_35_2: value  <=  10;
            Y_COORD_8_36_0: value  <=  4;
            Y_COORD_8_36_1: value  <=  5;
            Y_COORD_8_37_0: value  <=  3;
            Y_COORD_8_37_1: value  <=  3;
            Y_COORD_8_38_0: value  <=  6;
            Y_COORD_8_38_1: value  <=  7;
            Y_COORD_8_39_0: value  <=  3;
            Y_COORD_8_39_1: value  <=  3;
            Y_COORD_8_40_0: value  <=  1;
            Y_COORD_8_40_1: value  <=  1;
            Y_COORD_8_40_2: value  <=  6;
            Y_COORD_8_41_0: value  <=  7;
            Y_COORD_8_41_1: value  <=  7;
            Y_COORD_8_42_0: value  <=  7;
            Y_COORD_8_42_1: value  <=  7;
            Y_COORD_8_43_0: value  <=  12;
            Y_COORD_8_43_1: value  <=  13;
            Y_COORD_8_44_0: value  <=  8;
            Y_COORD_8_44_1: value  <=  8;
            Y_COORD_8_45_0: value  <=  4;
            Y_COORD_8_45_1: value  <=  10;
            Y_COORD_8_46_0: value  <=  5;
            Y_COORD_8_46_1: value  <=  5;
            Y_COORD_8_46_2: value  <=  11;
            Y_COORD_8_47_0: value  <=  14;
            Y_COORD_8_47_1: value  <=  15;
            Y_COORD_8_48_0: value  <=  12;
            Y_COORD_8_48_1: value  <=  13;
            Y_COORD_8_49_0: value  <=  2;
            Y_COORD_8_49_1: value  <=  2;
            Y_COORD_8_49_2: value  <=  3;
            Y_COORD_8_50_0: value  <=  1;
            Y_COORD_8_50_1: value  <=  1;
            Y_COORD_8_51_0: value  <=  0;
            Y_COORD_8_51_1: value  <=  0;
            Y_COORD_8_52_0: value  <=  7;
            Y_COORD_8_52_1: value  <=  7;
            Y_COORD_8_53_0: value  <=  1;
            Y_COORD_8_53_1: value  <=  6;
            Y_COORD_8_54_0: value  <=  1;
            Y_COORD_8_54_1: value  <=  1;
            Y_COORD_8_55_0: value  <=  3;
            Y_COORD_8_55_1: value  <=  5;
            Y_COORD_9_0_0: value  <=  3;
            Y_COORD_9_0_1: value  <=  6;
            Y_COORD_9_1_0: value  <=  7;
            Y_COORD_9_1_1: value  <=  7;
            Y_COORD_9_2_0: value  <=  4;
            Y_COORD_9_2_1: value  <=  9;
            Y_COORD_9_3_0: value  <=  4;
            Y_COORD_9_3_1: value  <=  12;
            Y_COORD_9_4_0: value  <=  15;
            Y_COORD_9_4_1: value  <=  17;
            Y_COORD_9_5_0: value  <=  2;
            Y_COORD_9_5_1: value  <=  2;
            Y_COORD_9_6_0: value  <=  3;
            Y_COORD_9_6_1: value  <=  4;
            Y_COORD_9_7_0: value  <=  6;
            Y_COORD_9_7_1: value  <=  9;
            Y_COORD_9_8_0: value  <=  11;
            Y_COORD_9_8_1: value  <=  12;
            Y_COORD_9_9_0: value  <=  2;
            Y_COORD_9_9_1: value  <=  2;
            Y_COORD_9_9_2: value  <=  5;
            Y_COORD_9_10_0: value  <=  2;
            Y_COORD_9_10_1: value  <=  2;
            Y_COORD_9_10_2: value  <=  7;
            Y_COORD_9_11_0: value  <=  10;
            Y_COORD_9_11_1: value  <=  12;
            Y_COORD_9_12_0: value  <=  10;
            Y_COORD_9_12_1: value  <=  12;
            Y_COORD_9_13_0: value  <=  5;
            Y_COORD_9_13_1: value  <=  5;
            Y_COORD_9_14_0: value  <=  6;
            Y_COORD_9_14_1: value  <=  10;
            Y_COORD_9_15_0: value  <=  11;
            Y_COORD_9_15_1: value  <=  14;
            Y_COORD_9_16_0: value  <=  13;
            Y_COORD_9_16_1: value  <=  13;
            Y_COORD_9_16_2: value  <=  16;
            Y_COORD_9_17_0: value  <=  0;
            Y_COORD_9_17_1: value  <=  0;
            Y_COORD_9_17_2: value  <=  6;
            Y_COORD_9_18_0: value  <=  0;
            Y_COORD_9_18_1: value  <=  1;
            Y_COORD_9_19_0: value  <=  12;
            Y_COORD_9_19_1: value  <=  13;
            Y_COORD_9_20_0: value  <=  12;
            Y_COORD_9_20_1: value  <=  13;
            Y_COORD_9_21_0: value  <=  11;
            Y_COORD_9_21_1: value  <=  12;
            Y_COORD_9_22_0: value  <=  3;
            Y_COORD_9_22_1: value  <=  3;
            Y_COORD_9_23_0: value  <=  7;
            Y_COORD_9_23_1: value  <=  9;
            Y_COORD_9_24_0: value  <=  2;
            Y_COORD_9_24_1: value  <=  2;
            Y_COORD_9_25_0: value  <=  4;
            Y_COORD_9_25_1: value  <=  5;
            Y_COORD_9_26_0: value  <=  4;
            Y_COORD_9_26_1: value  <=  5;
            Y_COORD_9_27_0: value  <=  3;
            Y_COORD_9_27_1: value  <=  4;
            Y_COORD_9_28_0: value  <=  5;
            Y_COORD_9_28_1: value  <=  6;
            Y_COORD_9_29_0: value  <=  7;
            Y_COORD_9_29_1: value  <=  9;
            Y_COORD_9_30_0: value  <=  7;
            Y_COORD_9_30_1: value  <=  9;
            Y_COORD_9_31_0: value  <=  2;
            Y_COORD_9_31_1: value  <=  5;
            Y_COORD_9_32_0: value  <=  4;
            Y_COORD_9_32_1: value  <=  6;
            Y_COORD_9_33_0: value  <=  5;
            Y_COORD_9_33_1: value  <=  5;
            Y_COORD_9_34_0: value  <=  5;
            Y_COORD_9_34_1: value  <=  5;
            Y_COORD_9_35_0: value  <=  1;
            Y_COORD_9_35_1: value  <=  3;
            Y_COORD_9_36_0: value  <=  2;
            Y_COORD_9_36_1: value  <=  4;
            Y_COORD_9_37_0: value  <=  6;
            Y_COORD_9_37_1: value  <=  7;
            Y_COORD_9_38_0: value  <=  1;
            Y_COORD_9_38_1: value  <=  4;
            Y_COORD_9_39_0: value  <=  0;
            Y_COORD_9_39_1: value  <=  0;
            Y_COORD_9_40_0: value  <=  10;
            Y_COORD_9_40_1: value  <=  11;
            Y_COORD_9_41_0: value  <=  4;
            Y_COORD_9_41_1: value  <=  9;
            Y_COORD_9_42_0: value  <=  1;
            Y_COORD_9_42_1: value  <=  1;
            Y_COORD_9_43_0: value  <=  11;
            Y_COORD_9_43_1: value  <=  11;
            Y_COORD_9_44_0: value  <=  11;
            Y_COORD_9_44_1: value  <=  11;
            Y_COORD_9_45_0: value  <=  8;
            Y_COORD_9_45_1: value  <=  8;
            Y_COORD_9_46_0: value  <=  0;
            Y_COORD_9_46_1: value  <=  0;
            Y_COORD_9_47_0: value  <=  4;
            Y_COORD_9_47_1: value  <=  4;
            Y_COORD_9_48_0: value  <=  12;
            Y_COORD_9_48_1: value  <=  16;
            Y_COORD_9_49_0: value  <=  14;
            Y_COORD_9_49_1: value  <=  15;
            Y_COORD_9_50_0: value  <=  14;
            Y_COORD_9_50_1: value  <=  15;
            Y_COORD_9_51_0: value  <=  4;
            Y_COORD_9_51_1: value  <=  4;
            Y_COORD_9_52_0: value  <=  15;
            Y_COORD_9_52_1: value  <=  15;
            Y_COORD_9_52_2: value  <=  17;
            Y_COORD_9_53_0: value  <=  2;
            Y_COORD_9_53_1: value  <=  2;
            Y_COORD_9_53_2: value  <=  4;
            Y_COORD_9_54_0: value  <=  8;
            Y_COORD_9_54_1: value  <=  8;
            Y_COORD_9_55_0: value  <=  7;
            Y_COORD_9_55_1: value  <=  7;
            Y_COORD_9_56_0: value  <=  7;
            Y_COORD_9_56_1: value  <=  7;
            Y_COORD_9_57_0: value  <=  7;
            Y_COORD_9_57_1: value  <=  7;
            Y_COORD_9_57_2: value  <=  9;
            Y_COORD_9_58_0: value  <=  13;
            Y_COORD_9_58_1: value  <=  14;
            Y_COORD_9_59_0: value  <=  7;
            Y_COORD_9_59_1: value  <=  7;
            Y_COORD_9_59_2: value  <=  9;
            Y_COORD_9_60_0: value  <=  7;
            Y_COORD_9_60_1: value  <=  7;
            Y_COORD_9_60_2: value  <=  9;
            Y_COORD_9_61_0: value  <=  6;
            Y_COORD_9_61_1: value  <=  12;
            Y_COORD_9_62_0: value  <=  5;
            Y_COORD_9_62_1: value  <=  5;
            Y_COORD_9_63_0: value  <=  12;
            Y_COORD_9_63_1: value  <=  13;
            Y_COORD_9_64_0: value  <=  12;
            Y_COORD_9_64_1: value  <=  13;
            Y_COORD_9_65_0: value  <=  12;
            Y_COORD_9_65_1: value  <=  13;
            Y_COORD_9_66_0: value  <=  2;
            Y_COORD_9_66_1: value  <=  2;
            Y_COORD_9_66_2: value  <=  4;
            Y_COORD_9_67_0: value  <=  5;
            Y_COORD_9_67_1: value  <=  6;
            Y_COORD_9_68_0: value  <=  6;
            Y_COORD_9_68_1: value  <=  12;
            Y_COORD_9_69_0: value  <=  13;
            Y_COORD_9_69_1: value  <=  13;
            Y_COORD_9_70_0: value  <=  6;
            Y_COORD_9_70_1: value  <=  12;
            Y_COORD_10_0_0: value  <=  2;
            Y_COORD_10_0_1: value  <=  2;
            Y_COORD_10_1_0: value  <=  5;
            Y_COORD_10_1_1: value  <=  5;
            Y_COORD_10_1_2: value  <=  10;
            Y_COORD_10_2_0: value  <=  5;
            Y_COORD_10_2_1: value  <=  5;
            Y_COORD_10_2_2: value  <=  11;
            Y_COORD_10_3_0: value  <=  7;
            Y_COORD_10_3_1: value  <=  9;
            Y_COORD_10_4_0: value  <=  2;
            Y_COORD_10_4_1: value  <=  3;
            Y_COORD_10_5_0: value  <=  18;
            Y_COORD_10_5_1: value  <=  18;
            Y_COORD_10_6_0: value  <=  4;
            Y_COORD_10_6_1: value  <=  12;
            Y_COORD_10_7_0: value  <=  6;
            Y_COORD_10_7_1: value  <=  10;
            Y_COORD_10_8_0: value  <=  3;
            Y_COORD_10_8_1: value  <=  3;
            Y_COORD_10_9_0: value  <=  15;
            Y_COORD_10_9_1: value  <=  17;
            Y_COORD_10_10_0: value  <=  5;
            Y_COORD_10_10_1: value  <=  9;
            Y_COORD_10_11_0: value  <=  1;
            Y_COORD_10_11_1: value  <=  7;
            Y_COORD_10_12_0: value  <=  6;
            Y_COORD_10_12_1: value  <=  6;
            Y_COORD_10_13_0: value  <=  4;
            Y_COORD_10_13_1: value  <=  6;
            Y_COORD_10_14_0: value  <=  3;
            Y_COORD_10_14_1: value  <=  4;
            Y_COORD_10_15_0: value  <=  11;
            Y_COORD_10_15_1: value  <=  12;
            Y_COORD_10_16_0: value  <=  16;
            Y_COORD_10_16_1: value  <=  17;
            Y_COORD_10_17_0: value  <=  13;
            Y_COORD_10_17_1: value  <=  13;
            Y_COORD_10_17_2: value  <=  16;
            Y_COORD_10_18_0: value  <=  0;
            Y_COORD_10_18_1: value  <=  0;
            Y_COORD_10_19_0: value  <=  15;
            Y_COORD_10_19_1: value  <=  16;
            Y_COORD_10_20_0: value  <=  4;
            Y_COORD_10_20_1: value  <=  6;
            Y_COORD_10_21_0: value  <=  6;
            Y_COORD_10_21_1: value  <=  6;
            Y_COORD_10_22_0: value  <=  6;
            Y_COORD_10_22_1: value  <=  6;
            Y_COORD_10_23_0: value  <=  7;
            Y_COORD_10_23_1: value  <=  7;
            Y_COORD_10_24_0: value  <=  12;
            Y_COORD_10_24_1: value  <=  14;
            Y_COORD_10_25_0: value  <=  12;
            Y_COORD_10_25_1: value  <=  14;
            Y_COORD_10_26_0: value  <=  0;
            Y_COORD_10_26_1: value  <=  1;
            Y_COORD_10_27_0: value  <=  0;
            Y_COORD_10_27_1: value  <=  0;
            Y_COORD_10_28_0: value  <=  3;
            Y_COORD_10_28_1: value  <=  3;
            Y_COORD_10_29_0: value  <=  0;
            Y_COORD_10_29_1: value  <=  0;
            Y_COORD_10_30_0: value  <=  3;
            Y_COORD_10_30_1: value  <=  8;
            Y_COORD_10_31_0: value  <=  0;
            Y_COORD_10_31_1: value  <=  0;
            Y_COORD_10_32_0: value  <=  0;
            Y_COORD_10_32_1: value  <=  0;
            Y_COORD_10_33_0: value  <=  15;
            Y_COORD_10_33_1: value  <=  16;
            Y_COORD_10_34_0: value  <=  2;
            Y_COORD_10_34_1: value  <=  2;
            Y_COORD_10_35_0: value  <=  1;
            Y_COORD_10_35_1: value  <=  1;
            Y_COORD_10_35_2: value  <=  3;
            Y_COORD_10_36_0: value  <=  12;
            Y_COORD_10_36_1: value  <=  13;
            Y_COORD_10_37_0: value  <=  2;
            Y_COORD_10_37_1: value  <=  2;
            Y_COORD_10_37_2: value  <=  5;
            Y_COORD_10_38_0: value  <=  7;
            Y_COORD_10_38_1: value  <=  7;
            Y_COORD_10_39_0: value  <=  7;
            Y_COORD_10_39_1: value  <=  7;
            Y_COORD_10_40_0: value  <=  5;
            Y_COORD_10_40_1: value  <=  5;
            Y_COORD_10_41_0: value  <=  15;
            Y_COORD_10_41_1: value  <=  16;
            Y_COORD_10_42_0: value  <=  18;
            Y_COORD_10_42_1: value  <=  18;
            Y_COORD_10_43_0: value  <=  13;
            Y_COORD_10_43_1: value  <=  14;
            Y_COORD_10_44_0: value  <=  13;
            Y_COORD_10_44_1: value  <=  14;
            Y_COORD_10_45_0: value  <=  15;
            Y_COORD_10_45_1: value  <=  16;
            Y_COORD_10_46_0: value  <=  15;
            Y_COORD_10_46_1: value  <=  17;
            Y_COORD_10_47_0: value  <=  3;
            Y_COORD_10_47_1: value  <=  3;
            Y_COORD_10_48_0: value  <=  14;
            Y_COORD_10_48_1: value  <=  15;
            Y_COORD_10_49_0: value  <=  14;
            Y_COORD_10_49_1: value  <=  16;
            Y_COORD_10_50_0: value  <=  3;
            Y_COORD_10_50_1: value  <=  6;
            Y_COORD_10_51_0: value  <=  11;
            Y_COORD_10_51_1: value  <=  14;
            Y_COORD_10_52_0: value  <=  10;
            Y_COORD_10_52_1: value  <=  10;
            Y_COORD_10_53_0: value  <=  9;
            Y_COORD_10_53_1: value  <=  9;
            Y_COORD_10_54_0: value  <=  3;
            Y_COORD_10_54_1: value  <=  3;
            Y_COORD_10_55_0: value  <=  7;
            Y_COORD_10_55_1: value  <=  7;
            Y_COORD_10_56_0: value  <=  12;
            Y_COORD_10_56_1: value  <=  13;
            Y_COORD_10_57_0: value  <=  8;
            Y_COORD_10_57_1: value  <=  12;
            Y_COORD_10_58_0: value  <=  14;
            Y_COORD_10_58_1: value  <=  14;
            Y_COORD_10_58_2: value  <=  17;
            Y_COORD_10_59_0: value  <=  15;
            Y_COORD_10_59_1: value  <=  16;
            Y_COORD_10_60_0: value  <=  15;
            Y_COORD_10_60_1: value  <=  16;
            Y_COORD_10_61_0: value  <=  12;
            Y_COORD_10_61_1: value  <=  13;
            Y_COORD_10_62_0: value  <=  7;
            Y_COORD_10_62_1: value  <=  7;
            Y_COORD_10_63_0: value  <=  6;
            Y_COORD_10_63_1: value  <=  6;
            Y_COORD_10_64_0: value  <=  7;
            Y_COORD_10_64_1: value  <=  7;
            Y_COORD_10_65_0: value  <=  7;
            Y_COORD_10_65_1: value  <=  7;
            Y_COORD_10_66_0: value  <=  7;
            Y_COORD_10_66_1: value  <=  7;
            Y_COORD_10_67_0: value  <=  1;
            Y_COORD_10_67_1: value  <=  1;
            Y_COORD_10_68_0: value  <=  2;
            Y_COORD_10_68_1: value  <=  2;
            Y_COORD_10_69_0: value  <=  14;
            Y_COORD_10_69_1: value  <=  14;
            Y_COORD_10_70_0: value  <=  8;
            Y_COORD_10_70_1: value  <=  9;
            Y_COORD_10_71_0: value  <=  7;
            Y_COORD_10_71_1: value  <=  8;
            Y_COORD_10_72_0: value  <=  6;
            Y_COORD_10_72_1: value  <=  6;
            Y_COORD_10_72_2: value  <=  7;
            Y_COORD_10_73_0: value  <=  11;
            Y_COORD_10_73_1: value  <=  11;
            Y_COORD_10_73_2: value  <=  13;
            Y_COORD_10_74_0: value  <=  6;
            Y_COORD_10_74_1: value  <=  6;
            Y_COORD_10_74_2: value  <=  7;
            Y_COORD_10_75_0: value  <=  15;
            Y_COORD_10_75_1: value  <=  16;
            Y_COORD_10_76_0: value  <=  14;
            Y_COORD_10_76_1: value  <=  15;
            Y_COORD_10_77_0: value  <=  14;
            Y_COORD_10_77_1: value  <=  15;
            Y_COORD_10_78_0: value  <=  7;
            Y_COORD_10_78_1: value  <=  8;
            Y_COORD_10_79_0: value  <=  10;
            Y_COORD_10_79_1: value  <=  11;
            Y_COORD_11_0_0: value  <=  4;
            Y_COORD_11_0_1: value  <=  6;
            Y_COORD_11_1_0: value  <=  7;
            Y_COORD_11_1_1: value  <=  7;
            Y_COORD_11_1_2: value  <=  9;
            Y_COORD_11_2_0: value  <=  7;
            Y_COORD_11_2_1: value  <=  9;
            Y_COORD_11_3_0: value  <=  15;
            Y_COORD_11_3_1: value  <=  15;
            Y_COORD_11_3_2: value  <=  17;
            Y_COORD_11_4_0: value  <=  8;
            Y_COORD_11_4_1: value  <=  9;
            Y_COORD_11_5_0: value  <=  1;
            Y_COORD_11_5_1: value  <=  1;
            Y_COORD_11_6_0: value  <=  15;
            Y_COORD_11_6_1: value  <=  15;
            Y_COORD_11_6_2: value  <=  17;
            Y_COORD_11_7_0: value  <=  5;
            Y_COORD_11_7_1: value  <=  5;
            Y_COORD_11_8_0: value  <=  6;
            Y_COORD_11_8_1: value  <=  6;
            Y_COORD_11_9_0: value  <=  9;
            Y_COORD_11_9_1: value  <=  10;
            Y_COORD_11_10_0: value  <=  15;
            Y_COORD_11_10_1: value  <=  16;
            Y_COORD_11_11_0: value  <=  10;
            Y_COORD_11_11_1: value  <=  10;
            Y_COORD_11_12_0: value  <=  9;
            Y_COORD_11_12_1: value  <=  14;
            Y_COORD_11_13_0: value  <=  11;
            Y_COORD_11_13_1: value  <=  11;
            Y_COORD_11_14_0: value  <=  11;
            Y_COORD_11_14_1: value  <=  11;
            Y_COORD_11_15_0: value  <=  3;
            Y_COORD_11_15_1: value  <=  3;
            Y_COORD_11_16_0: value  <=  3;
            Y_COORD_11_16_1: value  <=  3;
            Y_COORD_11_17_0: value  <=  5;
            Y_COORD_11_17_1: value  <=  5;
            Y_COORD_11_18_0: value  <=  5;
            Y_COORD_11_18_1: value  <=  11;
            Y_COORD_11_19_0: value  <=  11;
            Y_COORD_11_19_1: value  <=  12;
            Y_COORD_11_20_0: value  <=  1;
            Y_COORD_11_20_1: value  <=  1;
            Y_COORD_11_21_0: value  <=  3;
            Y_COORD_11_21_1: value  <=  5;
            Y_COORD_11_22_0: value  <=  3;
            Y_COORD_11_22_1: value  <=  5;
            Y_COORD_11_23_0: value  <=  12;
            Y_COORD_11_23_1: value  <=  13;
            Y_COORD_11_24_0: value  <=  13;
            Y_COORD_11_24_1: value  <=  14;
            Y_COORD_11_25_0: value  <=  0;
            Y_COORD_11_25_1: value  <=  2;
            Y_COORD_11_26_0: value  <=  0;
            Y_COORD_11_26_1: value  <=  2;
            Y_COORD_11_27_0: value  <=  14;
            Y_COORD_11_27_1: value  <=  15;
            Y_COORD_11_28_0: value  <=  4;
            Y_COORD_11_28_1: value  <=  4;
            Y_COORD_11_29_0: value  <=  5;
            Y_COORD_11_29_1: value  <=  7;
            Y_COORD_11_30_0: value  <=  4;
            Y_COORD_11_30_1: value  <=  4;
            Y_COORD_11_31_0: value  <=  14;
            Y_COORD_11_31_1: value  <=  14;
            Y_COORD_11_31_2: value  <=  16;
            Y_COORD_11_32_0: value  <=  15;
            Y_COORD_11_32_1: value  <=  15;
            Y_COORD_11_32_2: value  <=  16;
            Y_COORD_11_33_0: value  <=  15;
            Y_COORD_11_33_1: value  <=  16;
            Y_COORD_11_34_0: value  <=  12;
            Y_COORD_11_34_1: value  <=  16;
            Y_COORD_11_35_0: value  <=  7;
            Y_COORD_11_35_1: value  <=  8;
            Y_COORD_11_36_0: value  <=  2;
            Y_COORD_11_36_1: value  <=  3;
            Y_COORD_11_37_0: value  <=  6;
            Y_COORD_11_37_1: value  <=  6;
            Y_COORD_11_38_0: value  <=  5;
            Y_COORD_11_38_1: value  <=  5;
            Y_COORD_11_39_0: value  <=  6;
            Y_COORD_11_39_1: value  <=  6;
            Y_COORD_11_40_0: value  <=  13;
            Y_COORD_11_40_1: value  <=  14;
            Y_COORD_11_41_0: value  <=  4;
            Y_COORD_11_41_1: value  <=  4;
            Y_COORD_11_42_0: value  <=  4;
            Y_COORD_11_42_1: value  <=  4;
            Y_COORD_11_43_0: value  <=  11;
            Y_COORD_11_43_1: value  <=  12;
            Y_COORD_11_44_0: value  <=  2;
            Y_COORD_11_44_1: value  <=  2;
            Y_COORD_11_45_0: value  <=  6;
            Y_COORD_11_45_1: value  <=  6;
            Y_COORD_11_46_0: value  <=  6;
            Y_COORD_11_46_1: value  <=  6;
            Y_COORD_11_46_2: value  <=  10;
            Y_COORD_11_47_0: value  <=  0;
            Y_COORD_11_47_1: value  <=  0;
            Y_COORD_11_48_0: value  <=  4;
            Y_COORD_11_48_1: value  <=  4;
            Y_COORD_11_48_2: value  <=  10;
            Y_COORD_11_49_0: value  <=  4;
            Y_COORD_11_49_1: value  <=  5;
            Y_COORD_11_50_0: value  <=  11;
            Y_COORD_11_50_1: value  <=  12;
            Y_COORD_11_51_0: value  <=  7;
            Y_COORD_11_51_1: value  <=  7;
            Y_COORD_11_52_0: value  <=  7;
            Y_COORD_11_52_1: value  <=  7;
            Y_COORD_11_53_0: value  <=  17;
            Y_COORD_11_53_1: value  <=  17;
            Y_COORD_11_54_0: value  <=  6;
            Y_COORD_11_54_1: value  <=  7;
            Y_COORD_11_55_0: value  <=  0;
            Y_COORD_11_55_1: value  <=  0;
            Y_COORD_11_56_0: value  <=  6;
            Y_COORD_11_56_1: value  <=  6;
            Y_COORD_11_56_2: value  <=  7;
            Y_COORD_11_57_0: value  <=  16;
            Y_COORD_11_57_1: value  <=  17;
            Y_COORD_11_58_0: value  <=  12;
            Y_COORD_11_58_1: value  <=  13;
            Y_COORD_11_59_0: value  <=  12;
            Y_COORD_11_59_1: value  <=  13;
            Y_COORD_11_60_0: value  <=  11;
            Y_COORD_11_60_1: value  <=  11;
            Y_COORD_11_60_2: value  <=  13;
            Y_COORD_11_61_0: value  <=  4;
            Y_COORD_11_61_1: value  <=  5;
            Y_COORD_11_62_0: value  <=  4;
            Y_COORD_11_62_1: value  <=  5;
            Y_COORD_11_63_0: value  <=  16;
            Y_COORD_11_63_1: value  <=  17;
            Y_COORD_11_64_0: value  <=  4;
            Y_COORD_11_64_1: value  <=  5;
            Y_COORD_11_65_0: value  <=  0;
            Y_COORD_11_65_1: value  <=  1;
            Y_COORD_11_66_0: value  <=  9;
            Y_COORD_11_66_1: value  <=  10;
            Y_COORD_11_67_0: value  <=  8;
            Y_COORD_11_67_1: value  <=  9;
            Y_COORD_11_68_0: value  <=  13;
            Y_COORD_11_68_1: value  <=  13;
            Y_COORD_11_69_0: value  <=  14;
            Y_COORD_11_69_1: value  <=  15;
            Y_COORD_11_70_0: value  <=  18;
            Y_COORD_11_70_1: value  <=  18;
            Y_COORD_11_71_0: value  <=  14;
            Y_COORD_11_71_1: value  <=  15;
            Y_COORD_11_72_0: value  <=  14;
            Y_COORD_11_72_1: value  <=  15;
            Y_COORD_11_73_0: value  <=  14;
            Y_COORD_11_73_1: value  <=  15;
            Y_COORD_11_74_0: value  <=  14;
            Y_COORD_11_74_1: value  <=  15;
            Y_COORD_11_75_0: value  <=  6;
            Y_COORD_11_75_1: value  <=  6;
            Y_COORD_11_76_0: value  <=  6;
            Y_COORD_11_76_1: value  <=  6;
            Y_COORD_11_77_0: value  <=  5;
            Y_COORD_11_77_1: value  <=  6;
            Y_COORD_11_78_0: value  <=  16;
            Y_COORD_11_78_1: value  <=  16;
            Y_COORD_11_79_0: value  <=  12;
            Y_COORD_11_79_1: value  <=  13;
            Y_COORD_11_80_0: value  <=  0;
            Y_COORD_11_80_1: value  <=  0;
            Y_COORD_11_81_0: value  <=  0;
            Y_COORD_11_81_1: value  <=  9;
            Y_COORD_11_82_0: value  <=  1;
            Y_COORD_11_82_1: value  <=  8;
            Y_COORD_11_83_0: value  <=  9;
            Y_COORD_11_83_1: value  <=  9;
            Y_COORD_11_84_0: value  <=  12;
            Y_COORD_11_84_1: value  <=  13;
            Y_COORD_11_85_0: value  <=  15;
            Y_COORD_11_85_1: value  <=  16;
            Y_COORD_11_86_0: value  <=  3;
            Y_COORD_11_86_1: value  <=  3;
            Y_COORD_11_86_2: value  <=  10;
            Y_COORD_11_87_0: value  <=  2;
            Y_COORD_11_87_1: value  <=  2;
            Y_COORD_11_87_2: value  <=  11;
            Y_COORD_11_88_0: value  <=  15;
            Y_COORD_11_88_1: value  <=  16;
            Y_COORD_11_89_0: value  <=  2;
            Y_COORD_11_89_1: value  <=  2;
            Y_COORD_11_89_2: value  <=  11;
            Y_COORD_11_90_0: value  <=  1;
            Y_COORD_11_90_1: value  <=  2;
            Y_COORD_11_91_0: value  <=  11;
            Y_COORD_11_91_1: value  <=  12;
            Y_COORD_11_92_0: value  <=  11;
            Y_COORD_11_92_1: value  <=  14;
            Y_COORD_11_93_0: value  <=  0;
            Y_COORD_11_93_1: value  <=  0;
            Y_COORD_11_94_0: value  <=  0;
            Y_COORD_11_94_1: value  <=  0;
            Y_COORD_11_95_0: value  <=  3;
            Y_COORD_11_95_1: value  <=  3;
            Y_COORD_11_96_0: value  <=  3;
            Y_COORD_11_96_1: value  <=  3;
            Y_COORD_11_97_0: value  <=  8;
            Y_COORD_11_97_1: value  <=  12;
            Y_COORD_11_98_0: value  <=  0;
            Y_COORD_11_98_1: value  <=  0;
            Y_COORD_11_99_0: value  <=  0;
            Y_COORD_11_99_1: value  <=  0;
            Y_COORD_11_100_0: value  <=  3;
            Y_COORD_11_100_1: value  <=  4;
            Y_COORD_11_101_0: value  <=  5;
            Y_COORD_11_101_1: value  <=  5;
            Y_COORD_11_101_2: value  <=  9;
            Y_COORD_11_102_0: value  <=  7;
            Y_COORD_11_102_1: value  <=  7;
            Y_COORD_11_102_2: value  <=  9;
            Y_COORD_12_0_0: value  <=  1;
            Y_COORD_12_0_1: value  <=  1;
            Y_COORD_12_1_0: value  <=  7;
            Y_COORD_12_1_1: value  <=  7;
            Y_COORD_12_1_2: value  <=  9;
            Y_COORD_12_2_0: value  <=  6;
            Y_COORD_12_2_1: value  <=  9;
            Y_COORD_12_3_0: value  <=  16;
            Y_COORD_12_3_1: value  <=  16;
            Y_COORD_12_3_2: value  <=  18;
            Y_COORD_12_4_0: value  <=  4;
            Y_COORD_12_4_1: value  <=  10;
            Y_COORD_12_5_0: value  <=  1;
            Y_COORD_12_5_1: value  <=  1;
            Y_COORD_12_6_0: value  <=  12;
            Y_COORD_12_6_1: value  <=  12;
            Y_COORD_12_7_0: value  <=  8;
            Y_COORD_12_7_1: value  <=  9;
            Y_COORD_12_8_0: value  <=  0;
            Y_COORD_12_8_1: value  <=  0;
            Y_COORD_12_9_0: value  <=  18;
            Y_COORD_12_9_1: value  <=  19;
            Y_COORD_12_10_0: value  <=  1;
            Y_COORD_12_10_1: value  <=  3;
            Y_COORD_12_11_0: value  <=  8;
            Y_COORD_12_11_1: value  <=  8;
            Y_COORD_12_12_0: value  <=  14;
            Y_COORD_12_12_1: value  <=  15;
            Y_COORD_12_13_0: value  <=  3;
            Y_COORD_12_13_1: value  <=  3;
            Y_COORD_12_14_0: value  <=  7;
            Y_COORD_12_14_1: value  <=  7;
            Y_COORD_12_15_0: value  <=  3;
            Y_COORD_12_15_1: value  <=  4;
            Y_COORD_12_16_0: value  <=  4;
            Y_COORD_12_16_1: value  <=  6;
            Y_COORD_12_17_0: value  <=  5;
            Y_COORD_12_17_1: value  <=  10;
            Y_COORD_12_18_0: value  <=  18;
            Y_COORD_12_18_1: value  <=  18;
            Y_COORD_12_19_0: value  <=  2;
            Y_COORD_12_19_1: value  <=  4;
            Y_COORD_12_20_0: value  <=  7;
            Y_COORD_12_20_1: value  <=  7;
            Y_COORD_12_21_0: value  <=  2;
            Y_COORD_12_21_1: value  <=  4;
            Y_COORD_12_22_0: value  <=  0;
            Y_COORD_12_22_1: value  <=  0;
            Y_COORD_12_23_0: value  <=  14;
            Y_COORD_12_23_1: value  <=  15;
            Y_COORD_12_24_0: value  <=  12;
            Y_COORD_12_24_1: value  <=  13;
            Y_COORD_12_25_0: value  <=  14;
            Y_COORD_12_25_1: value  <=  15;
            Y_COORD_12_26_0: value  <=  12;
            Y_COORD_12_26_1: value  <=  13;
            Y_COORD_12_27_0: value  <=  6;
            Y_COORD_12_27_1: value  <=  6;
            Y_COORD_12_28_0: value  <=  2;
            Y_COORD_12_28_1: value  <=  4;
            Y_COORD_12_29_0: value  <=  6;
            Y_COORD_12_29_1: value  <=  7;
            Y_COORD_12_30_0: value  <=  0;
            Y_COORD_12_30_1: value  <=  0;
            Y_COORD_12_31_0: value  <=  14;
            Y_COORD_12_31_1: value  <=  16;
            Y_COORD_12_32_0: value  <=  14;
            Y_COORD_12_32_1: value  <=  16;
            Y_COORD_12_33_0: value  <=  10;
            Y_COORD_12_33_1: value  <=  10;
            Y_COORD_12_33_2: value  <=  11;
            Y_COORD_12_34_0: value  <=  0;
            Y_COORD_12_34_1: value  <=  0;
            Y_COORD_12_35_0: value  <=  15;
            Y_COORD_12_35_1: value  <=  16;
            Y_COORD_12_36_0: value  <=  2;
            Y_COORD_12_36_1: value  <=  3;
            Y_COORD_12_37_0: value  <=  11;
            Y_COORD_12_37_1: value  <=  14;
            Y_COORD_12_38_0: value  <=  11;
            Y_COORD_12_38_1: value  <=  14;
            Y_COORD_12_39_0: value  <=  10;
            Y_COORD_12_39_1: value  <=  10;
            Y_COORD_12_39_2: value  <=  11;
            Y_COORD_12_40_0: value  <=  6;
            Y_COORD_12_40_1: value  <=  7;
            Y_COORD_12_41_0: value  <=  9;
            Y_COORD_12_41_1: value  <=  10;
            Y_COORD_12_42_0: value  <=  7;
            Y_COORD_12_42_1: value  <=  7;
            Y_COORD_12_43_0: value  <=  5;
            Y_COORD_12_43_1: value  <=  5;
            Y_COORD_12_44_0: value  <=  10;
            Y_COORD_12_44_1: value  <=  11;
            Y_COORD_12_45_0: value  <=  14;
            Y_COORD_12_45_1: value  <=  15;
            Y_COORD_12_46_0: value  <=  11;
            Y_COORD_12_46_1: value  <=  12;
            Y_COORD_12_47_0: value  <=  1;
            Y_COORD_12_47_1: value  <=  7;
            Y_COORD_12_48_0: value  <=  1;
            Y_COORD_12_48_1: value  <=  1;
            Y_COORD_12_48_2: value  <=  6;
            Y_COORD_12_49_0: value  <=  1;
            Y_COORD_12_49_1: value  <=  2;
            Y_COORD_12_50_0: value  <=  5;
            Y_COORD_12_50_1: value  <=  6;
            Y_COORD_12_51_0: value  <=  2;
            Y_COORD_12_51_1: value  <=  2;
            Y_COORD_12_52_0: value  <=  3;
            Y_COORD_12_52_1: value  <=  5;
            Y_COORD_12_53_0: value  <=  12;
            Y_COORD_12_53_1: value  <=  13;
            Y_COORD_12_54_0: value  <=  18;
            Y_COORD_12_54_1: value  <=  18;
            Y_COORD_12_55_0: value  <=  10;
            Y_COORD_12_55_1: value  <=  10;
            Y_COORD_12_55_2: value  <=  11;
            Y_COORD_12_56_0: value  <=  10;
            Y_COORD_12_56_1: value  <=  10;
            Y_COORD_12_56_2: value  <=  11;
            Y_COORD_12_57_0: value  <=  11;
            Y_COORD_12_57_1: value  <=  13;
            Y_COORD_12_58_0: value  <=  12;
            Y_COORD_12_58_1: value  <=  12;
            Y_COORD_12_59_0: value  <=  0;
            Y_COORD_12_59_1: value  <=  1;
            Y_COORD_12_60_0: value  <=  8;
            Y_COORD_12_60_1: value  <=  8;
            Y_COORD_12_61_0: value  <=  7;
            Y_COORD_12_61_1: value  <=  7;
            Y_COORD_12_61_2: value  <=  12;
            Y_COORD_12_62_0: value  <=  18;
            Y_COORD_12_62_1: value  <=  18;
            Y_COORD_12_62_2: value  <=  19;
            Y_COORD_12_63_0: value  <=  2;
            Y_COORD_12_63_1: value  <=  2;
            Y_COORD_12_64_0: value  <=  2;
            Y_COORD_12_64_1: value  <=  2;
            Y_COORD_12_65_0: value  <=  0;
            Y_COORD_12_65_1: value  <=  0;
            Y_COORD_12_66_0: value  <=  11;
            Y_COORD_12_66_1: value  <=  11;
            Y_COORD_12_67_0: value  <=  14;
            Y_COORD_12_67_1: value  <=  15;
            Y_COORD_12_68_0: value  <=  15;
            Y_COORD_12_68_1: value  <=  15;
            Y_COORD_12_68_2: value  <=  16;
            Y_COORD_12_69_0: value  <=  14;
            Y_COORD_12_69_1: value  <=  15;
            Y_COORD_12_70_0: value  <=  0;
            Y_COORD_12_70_1: value  <=  0;
            Y_COORD_12_71_0: value  <=  1;
            Y_COORD_12_71_1: value  <=  1;
            Y_COORD_12_72_0: value  <=  0;
            Y_COORD_12_72_1: value  <=  10;
            Y_COORD_12_73_0: value  <=  0;
            Y_COORD_12_73_1: value  <=  2;
            Y_COORD_12_74_0: value  <=  3;
            Y_COORD_12_74_1: value  <=  4;
            Y_COORD_12_75_0: value  <=  0;
            Y_COORD_12_75_1: value  <=  0;
            Y_COORD_12_76_0: value  <=  0;
            Y_COORD_12_76_1: value  <=  0;
            Y_COORD_12_77_0: value  <=  0;
            Y_COORD_12_77_1: value  <=  0;
            Y_COORD_12_78_0: value  <=  7;
            Y_COORD_12_78_1: value  <=  7;
            Y_COORD_12_79_0: value  <=  0;
            Y_COORD_12_79_1: value  <=  0;
            Y_COORD_12_80_0: value  <=  0;
            Y_COORD_12_80_1: value  <=  0;
            Y_COORD_12_81_0: value  <=  12;
            Y_COORD_12_81_1: value  <=  14;
            Y_COORD_12_82_0: value  <=  12;
            Y_COORD_12_82_1: value  <=  14;
            Y_COORD_12_83_0: value  <=  1;
            Y_COORD_12_83_1: value  <=  2;
            Y_COORD_12_84_0: value  <=  7;
            Y_COORD_12_84_1: value  <=  7;
            Y_COORD_12_84_2: value  <=  12;
            Y_COORD_12_85_0: value  <=  11;
            Y_COORD_12_85_1: value  <=  13;
            Y_COORD_12_86_0: value  <=  1;
            Y_COORD_12_86_1: value  <=  2;
            Y_COORD_12_87_0: value  <=  4;
            Y_COORD_12_87_1: value  <=  5;
            Y_COORD_12_88_0: value  <=  15;
            Y_COORD_12_88_1: value  <=  15;
            Y_COORD_12_89_0: value  <=  7;
            Y_COORD_12_89_1: value  <=  7;
            Y_COORD_12_90_0: value  <=  7;
            Y_COORD_12_90_1: value  <=  7;
            Y_COORD_12_91_0: value  <=  6;
            Y_COORD_12_91_1: value  <=  6;
            Y_COORD_12_92_0: value  <=  5;
            Y_COORD_12_92_1: value  <=  7;
            Y_COORD_12_93_0: value  <=  5;
            Y_COORD_12_93_1: value  <=  5;
            Y_COORD_12_94_0: value  <=  0;
            Y_COORD_12_94_1: value  <=  0;
            Y_COORD_12_95_0: value  <=  6;
            Y_COORD_12_95_1: value  <=  6;
            Y_COORD_12_96_0: value  <=  6;
            Y_COORD_12_96_1: value  <=  6;
            Y_COORD_12_97_0: value  <=  4;
            Y_COORD_12_97_1: value  <=  5;
            Y_COORD_12_98_0: value  <=  1;
            Y_COORD_12_98_1: value  <=  1;
            Y_COORD_12_99_0: value  <=  1;
            Y_COORD_12_99_1: value  <=  1;
            Y_COORD_12_99_2: value  <=  10;
            Y_COORD_12_100_0: value  <=  1;
            Y_COORD_12_100_1: value  <=  2;
            Y_COORD_12_101_0: value  <=  1;
            Y_COORD_12_101_1: value  <=  1;
            Y_COORD_12_101_2: value  <=  10;
            Y_COORD_12_102_0: value  <=  14;
            Y_COORD_12_102_1: value  <=  14;
            Y_COORD_12_102_2: value  <=  17;
            Y_COORD_12_103_0: value  <=  11;
            Y_COORD_12_103_1: value  <=  13;
            Y_COORD_12_104_0: value  <=  10;
            Y_COORD_12_104_1: value  <=  10;
            Y_COORD_12_104_2: value  <=  15;
            Y_COORD_12_105_0: value  <=  0;
            Y_COORD_12_105_1: value  <=  0;
            Y_COORD_12_106_0: value  <=  10;
            Y_COORD_12_106_1: value  <=  13;
            Y_COORD_12_107_0: value  <=  6;
            Y_COORD_12_107_1: value  <=  10;
            Y_COORD_12_108_0: value  <=  7;
            Y_COORD_12_108_1: value  <=  7;
            Y_COORD_12_108_2: value  <=  10;
            Y_COORD_12_109_0: value  <=  7;
            Y_COORD_12_109_1: value  <=  7;
            Y_COORD_12_110_0: value  <=  9;
            Y_COORD_12_110_1: value  <=  9;
            Y_COORD_13_0_0: value  <=  6;
            Y_COORD_13_0_1: value  <=  6;
            Y_COORD_13_1_0: value  <=  0;
            Y_COORD_13_1_1: value  <=  0;
            Y_COORD_13_2_0: value  <=  15;
            Y_COORD_13_2_1: value  <=  17;
            Y_COORD_13_3_0: value  <=  0;
            Y_COORD_13_3_1: value  <=  3;
            Y_COORD_13_4_0: value  <=  7;
            Y_COORD_13_4_1: value  <=  9;
            Y_COORD_13_5_0: value  <=  7;
            Y_COORD_13_5_1: value  <=  7;
            Y_COORD_13_5_2: value  <=  9;
            Y_COORD_13_6_0: value  <=  7;
            Y_COORD_13_6_1: value  <=  7;
            Y_COORD_13_6_2: value  <=  9;
            Y_COORD_13_7_0: value  <=  6;
            Y_COORD_13_7_1: value  <=  10;
            Y_COORD_13_8_0: value  <=  8;
            Y_COORD_13_8_1: value  <=  14;
            Y_COORD_13_9_0: value  <=  5;
            Y_COORD_13_9_1: value  <=  5;
            Y_COORD_13_9_2: value  <=  11;
            Y_COORD_13_10_0: value  <=  11;
            Y_COORD_13_10_1: value  <=  12;
            Y_COORD_13_11_0: value  <=  5;
            Y_COORD_13_11_1: value  <=  5;
            Y_COORD_13_12_0: value  <=  4;
            Y_COORD_13_12_1: value  <=  6;
            Y_COORD_13_13_0: value  <=  5;
            Y_COORD_13_13_1: value  <=  5;
            Y_COORD_13_14_0: value  <=  5;
            Y_COORD_13_14_1: value  <=  5;
            Y_COORD_13_15_0: value  <=  2;
            Y_COORD_13_15_1: value  <=  2;
            Y_COORD_13_16_0: value  <=  2;
            Y_COORD_13_16_1: value  <=  2;
            Y_COORD_13_17_0: value  <=  5;
            Y_COORD_13_17_1: value  <=  6;
            Y_COORD_13_18_0: value  <=  10;
            Y_COORD_13_18_1: value  <=  12;
            Y_COORD_13_19_0: value  <=  5;
            Y_COORD_13_19_1: value  <=  6;
            Y_COORD_13_20_0: value  <=  18;
            Y_COORD_13_20_1: value  <=  18;
            Y_COORD_13_21_0: value  <=  15;
            Y_COORD_13_21_1: value  <=  16;
            Y_COORD_13_22_0: value  <=  14;
            Y_COORD_13_22_1: value  <=  15;
            Y_COORD_13_23_0: value  <=  4;
            Y_COORD_13_23_1: value  <=  6;
            Y_COORD_13_24_0: value  <=  5;
            Y_COORD_13_24_1: value  <=  6;
            Y_COORD_13_25_0: value  <=  16;
            Y_COORD_13_25_1: value  <=  17;
            Y_COORD_13_26_0: value  <=  0;
            Y_COORD_13_26_1: value  <=  3;
            Y_COORD_13_27_0: value  <=  7;
            Y_COORD_13_27_1: value  <=  8;
            Y_COORD_13_28_0: value  <=  7;
            Y_COORD_13_28_1: value  <=  8;
            Y_COORD_13_29_0: value  <=  5;
            Y_COORD_13_29_1: value  <=  5;
            Y_COORD_13_30_0: value  <=  6;
            Y_COORD_13_30_1: value  <=  6;
            Y_COORD_13_31_0: value  <=  6;
            Y_COORD_13_31_1: value  <=  6;
            Y_COORD_13_31_2: value  <=  12;
            Y_COORD_13_32_0: value  <=  6;
            Y_COORD_13_32_1: value  <=  6;
            Y_COORD_13_32_2: value  <=  12;
            Y_COORD_13_33_0: value  <=  4;
            Y_COORD_13_33_1: value  <=  5;
            Y_COORD_13_34_0: value  <=  16;
            Y_COORD_13_34_1: value  <=  17;
            Y_COORD_13_35_0: value  <=  4;
            Y_COORD_13_35_1: value  <=  5;
            Y_COORD_13_36_0: value  <=  12;
            Y_COORD_13_36_1: value  <=  14;
            Y_COORD_13_37_0: value  <=  13;
            Y_COORD_13_37_1: value  <=  14;
            Y_COORD_13_38_0: value  <=  14;
            Y_COORD_13_38_1: value  <=  15;
            Y_COORD_13_39_0: value  <=  15;
            Y_COORD_13_39_1: value  <=  16;
            Y_COORD_13_40_0: value  <=  4;
            Y_COORD_13_40_1: value  <=  5;
            Y_COORD_13_41_0: value  <=  15;
            Y_COORD_13_41_1: value  <=  16;
            Y_COORD_13_42_0: value  <=  3;
            Y_COORD_13_42_1: value  <=  3;
            Y_COORD_13_43_0: value  <=  15;
            Y_COORD_13_43_1: value  <=  16;
            Y_COORD_13_44_0: value  <=  15;
            Y_COORD_13_44_1: value  <=  16;
            Y_COORD_13_45_0: value  <=  13;
            Y_COORD_13_45_1: value  <=  13;
            Y_COORD_13_45_2: value  <=  16;
            Y_COORD_13_46_0: value  <=  8;
            Y_COORD_13_46_1: value  <=  8;
            Y_COORD_13_47_0: value  <=  0;
            Y_COORD_13_47_1: value  <=  2;
            Y_COORD_13_48_0: value  <=  2;
            Y_COORD_13_48_1: value  <=  2;
            Y_COORD_13_48_2: value  <=  3;
            Y_COORD_13_49_0: value  <=  0;
            Y_COORD_13_49_1: value  <=  0;
            Y_COORD_13_50_0: value  <=  3;
            Y_COORD_13_50_1: value  <=  3;
            Y_COORD_13_51_0: value  <=  18;
            Y_COORD_13_51_1: value  <=  19;
            Y_COORD_13_52_0: value  <=  10;
            Y_COORD_13_52_1: value  <=  12;
            Y_COORD_13_53_0: value  <=  12;
            Y_COORD_13_53_1: value  <=  12;
            Y_COORD_13_53_2: value  <=  16;
            Y_COORD_13_54_0: value  <=  13;
            Y_COORD_13_54_1: value  <=  13;
            Y_COORD_13_54_2: value  <=  16;
            Y_COORD_13_55_0: value  <=  12;
            Y_COORD_13_55_1: value  <=  13;
            Y_COORD_13_56_0: value  <=  13;
            Y_COORD_13_56_1: value  <=  14;
            Y_COORD_13_57_0: value  <=  12;
            Y_COORD_13_57_1: value  <=  13;
            Y_COORD_13_58_0: value  <=  12;
            Y_COORD_13_58_1: value  <=  13;
            Y_COORD_13_59_0: value  <=  12;
            Y_COORD_13_59_1: value  <=  13;
            Y_COORD_13_60_0: value  <=  14;
            Y_COORD_13_60_1: value  <=  15;
            Y_COORD_13_61_0: value  <=  10;
            Y_COORD_13_61_1: value  <=  13;
            Y_COORD_13_62_0: value  <=  6;
            Y_COORD_13_62_1: value  <=  12;
            Y_COORD_13_63_0: value  <=  10;
            Y_COORD_13_63_1: value  <=  13;
            Y_COORD_13_64_0: value  <=  10;
            Y_COORD_13_64_1: value  <=  13;
            Y_COORD_13_65_0: value  <=  4;
            Y_COORD_13_65_1: value  <=  5;
            Y_COORD_13_66_0: value  <=  1;
            Y_COORD_13_66_1: value  <=  6;
            Y_COORD_13_67_0: value  <=  8;
            Y_COORD_13_67_1: value  <=  9;
            Y_COORD_13_68_0: value  <=  17;
            Y_COORD_13_68_1: value  <=  18;
            Y_COORD_13_69_0: value  <=  9;
            Y_COORD_13_69_1: value  <=  9;
            Y_COORD_13_70_0: value  <=  14;
            Y_COORD_13_70_1: value  <=  14;
            Y_COORD_13_70_2: value  <=  17;
            Y_COORD_13_71_0: value  <=  9;
            Y_COORD_13_71_1: value  <=  9;
            Y_COORD_13_72_0: value  <=  9;
            Y_COORD_13_72_1: value  <=  9;
            Y_COORD_13_73_0: value  <=  10;
            Y_COORD_13_73_1: value  <=  10;
            Y_COORD_13_74_0: value  <=  0;
            Y_COORD_13_74_1: value  <=  1;
            Y_COORD_13_75_0: value  <=  9;
            Y_COORD_13_75_1: value  <=  12;
            Y_COORD_13_76_0: value  <=  1;
            Y_COORD_13_76_1: value  <=  1;
            Y_COORD_13_77_0: value  <=  3;
            Y_COORD_13_77_1: value  <=  4;
            Y_COORD_13_78_0: value  <=  3;
            Y_COORD_13_78_1: value  <=  4;
            Y_COORD_13_79_0: value  <=  7;
            Y_COORD_13_79_1: value  <=  7;
            Y_COORD_13_80_0: value  <=  5;
            Y_COORD_13_80_1: value  <=  5;
            Y_COORD_13_81_0: value  <=  5;
            Y_COORD_13_81_1: value  <=  5;
            Y_COORD_13_82_0: value  <=  4;
            Y_COORD_13_82_1: value  <=  4;
            Y_COORD_13_82_2: value  <=  10;
            Y_COORD_13_83_0: value  <=  2;
            Y_COORD_13_83_1: value  <=  2;
            Y_COORD_13_84_0: value  <=  2;
            Y_COORD_13_84_1: value  <=  2;
            Y_COORD_13_85_0: value  <=  10;
            Y_COORD_13_85_1: value  <=  10;
            Y_COORD_13_86_0: value  <=  10;
            Y_COORD_13_86_1: value  <=  10;
            Y_COORD_13_87_0: value  <=  2;
            Y_COORD_13_87_1: value  <=  2;
            Y_COORD_13_88_0: value  <=  2;
            Y_COORD_13_88_1: value  <=  2;
            Y_COORD_13_89_0: value  <=  9;
            Y_COORD_13_89_1: value  <=  11;
            Y_COORD_13_90_0: value  <=  7;
            Y_COORD_13_90_1: value  <=  7;
            Y_COORD_13_91_0: value  <=  10;
            Y_COORD_13_91_1: value  <=  10;
            Y_COORD_13_91_2: value  <=  13;
            Y_COORD_13_92_0: value  <=  9;
            Y_COORD_13_92_1: value  <=  12;
            Y_COORD_13_93_0: value  <=  15;
            Y_COORD_13_93_1: value  <=  16;
            Y_COORD_13_94_0: value  <=  12;
            Y_COORD_13_94_1: value  <=  14;
            Y_COORD_13_95_0: value  <=  3;
            Y_COORD_13_95_1: value  <=  9;
            Y_COORD_13_96_0: value  <=  1;
            Y_COORD_13_96_1: value  <=  1;
            Y_COORD_13_96_2: value  <=  7;
            Y_COORD_13_97_0: value  <=  4;
            Y_COORD_13_97_1: value  <=  4;
            Y_COORD_13_97_2: value  <=  6;
            Y_COORD_13_98_0: value  <=  9;
            Y_COORD_13_98_1: value  <=  9;
            Y_COORD_13_98_2: value  <=  10;
            Y_COORD_13_99_0: value  <=  11;
            Y_COORD_13_99_1: value  <=  12;
            Y_COORD_13_100_0: value  <=  12;
            Y_COORD_13_100_1: value  <=  13;
            Y_COORD_13_101_0: value  <=  9;
            Y_COORD_13_101_1: value  <=  10;
            Y_COORD_14_0_0: value  <=  4;
            Y_COORD_14_0_1: value  <=  6;
            Y_COORD_14_1_0: value  <=  7;
            Y_COORD_14_1_1: value  <=  7;
            Y_COORD_14_1_2: value  <=  9;
            Y_COORD_14_2_0: value  <=  0;
            Y_COORD_14_2_1: value  <=  0;
            Y_COORD_14_3_0: value  <=  5;
            Y_COORD_14_3_1: value  <=  11;
            Y_COORD_14_4_0: value  <=  4;
            Y_COORD_14_4_1: value  <=  9;
            Y_COORD_14_5_0: value  <=  17;
            Y_COORD_14_5_1: value  <=  18;
            Y_COORD_14_6_0: value  <=  5;
            Y_COORD_14_6_1: value  <=  7;
            Y_COORD_14_7_0: value  <=  2;
            Y_COORD_14_7_1: value  <=  3;
            Y_COORD_14_8_0: value  <=  5;
            Y_COORD_14_8_1: value  <=  5;
            Y_COORD_14_9_0: value  <=  14;
            Y_COORD_14_9_1: value  <=  16;
            Y_COORD_14_10_0: value  <=  11;
            Y_COORD_14_10_1: value  <=  12;
            Y_COORD_14_11_0: value  <=  13;
            Y_COORD_14_11_1: value  <=  14;
            Y_COORD_14_12_0: value  <=  5;
            Y_COORD_14_12_1: value  <=  7;
            Y_COORD_14_13_0: value  <=  2;
            Y_COORD_14_13_1: value  <=  3;
            Y_COORD_14_14_0: value  <=  14;
            Y_COORD_14_14_1: value  <=  14;
            Y_COORD_14_14_2: value  <=  17;
            Y_COORD_14_15_0: value  <=  2;
            Y_COORD_14_15_1: value  <=  3;
            Y_COORD_14_16_0: value  <=  2;
            Y_COORD_14_16_1: value  <=  6;
            Y_COORD_14_17_0: value  <=  0;
            Y_COORD_14_17_1: value  <=  0;
            Y_COORD_14_17_2: value  <=  4;
            Y_COORD_14_18_0: value  <=  17;
            Y_COORD_14_18_1: value  <=  17;
            Y_COORD_14_19_0: value  <=  12;
            Y_COORD_14_19_1: value  <=  13;
            Y_COORD_14_20_0: value  <=  0;
            Y_COORD_14_20_1: value  <=  0;
            Y_COORD_14_20_2: value  <=  6;
            Y_COORD_14_21_0: value  <=  0;
            Y_COORD_14_21_1: value  <=  0;
            Y_COORD_14_21_2: value  <=  5;
            Y_COORD_14_22_0: value  <=  3;
            Y_COORD_14_22_1: value  <=  3;
            Y_COORD_14_22_2: value  <=  6;
            Y_COORD_14_23_0: value  <=  0;
            Y_COORD_14_23_1: value  <=  0;
            Y_COORD_14_23_2: value  <=  5;
            Y_COORD_14_24_0: value  <=  14;
            Y_COORD_14_24_1: value  <=  15;
            Y_COORD_14_25_0: value  <=  10;
            Y_COORD_14_25_1: value  <=  11;
            Y_COORD_14_26_0: value  <=  14;
            Y_COORD_14_26_1: value  <=  15;
            Y_COORD_14_27_0: value  <=  13;
            Y_COORD_14_27_1: value  <=  13;
            Y_COORD_14_27_2: value  <=  15;
            Y_COORD_14_28_0: value  <=  10;
            Y_COORD_14_28_1: value  <=  11;
            Y_COORD_14_29_0: value  <=  11;
            Y_COORD_14_29_1: value  <=  11;
            Y_COORD_14_30_0: value  <=  11;
            Y_COORD_14_30_1: value  <=  11;
            Y_COORD_14_31_0: value  <=  5;
            Y_COORD_14_31_1: value  <=  10;
            Y_COORD_14_32_0: value  <=  12;
            Y_COORD_14_32_1: value  <=  12;
            Y_COORD_14_33_0: value  <=  4;
            Y_COORD_14_33_1: value  <=  4;
            Y_COORD_14_33_2: value  <=  9;
            Y_COORD_14_34_0: value  <=  6;
            Y_COORD_14_34_1: value  <=  6;
            Y_COORD_14_35_0: value  <=  12;
            Y_COORD_14_35_1: value  <=  12;
            Y_COORD_14_35_2: value  <=  16;
            Y_COORD_14_36_0: value  <=  14;
            Y_COORD_14_36_1: value  <=  15;
            Y_COORD_14_37_0: value  <=  2;
            Y_COORD_14_37_1: value  <=  2;
            Y_COORD_14_38_0: value  <=  15;
            Y_COORD_14_38_1: value  <=  16;
            Y_COORD_14_39_0: value  <=  0;
            Y_COORD_14_39_1: value  <=  0;
            Y_COORD_14_40_0: value  <=  6;
            Y_COORD_14_40_1: value  <=  6;
            Y_COORD_14_41_0: value  <=  8;
            Y_COORD_14_41_1: value  <=  9;
            Y_COORD_14_42_0: value  <=  9;
            Y_COORD_14_42_1: value  <=  11;
            Y_COORD_14_43_0: value  <=  0;
            Y_COORD_14_43_1: value  <=  1;
            Y_COORD_14_44_0: value  <=  14;
            Y_COORD_14_44_1: value  <=  15;
            Y_COORD_14_45_0: value  <=  10;
            Y_COORD_14_45_1: value  <=  13;
            Y_COORD_14_46_0: value  <=  2;
            Y_COORD_14_46_1: value  <=  2;
            Y_COORD_14_47_0: value  <=  1;
            Y_COORD_14_47_1: value  <=  1;
            Y_COORD_14_47_2: value  <=  5;
            Y_COORD_14_48_0: value  <=  1;
            Y_COORD_14_48_1: value  <=  1;
            Y_COORD_14_48_2: value  <=  5;
            Y_COORD_14_49_0: value  <=  2;
            Y_COORD_14_49_1: value  <=  2;
            Y_COORD_14_49_2: value  <=  5;
            Y_COORD_14_50_0: value  <=  3;
            Y_COORD_14_50_1: value  <=  3;
            Y_COORD_14_51_0: value  <=  2;
            Y_COORD_14_51_1: value  <=  2;
            Y_COORD_14_51_2: value  <=  5;
            Y_COORD_14_52_0: value  <=  4;
            Y_COORD_14_52_1: value  <=  5;
            Y_COORD_14_53_0: value  <=  5;
            Y_COORD_14_53_1: value  <=  6;
            Y_COORD_14_54_0: value  <=  16;
            Y_COORD_14_54_1: value  <=  17;
            Y_COORD_14_55_0: value  <=  2;
            Y_COORD_14_55_1: value  <=  2;
            Y_COORD_14_55_2: value  <=  5;
            Y_COORD_14_56_0: value  <=  2;
            Y_COORD_14_56_1: value  <=  2;
            Y_COORD_14_56_2: value  <=  5;
            Y_COORD_14_57_0: value  <=  5;
            Y_COORD_14_57_1: value  <=  6;
            Y_COORD_14_58_0: value  <=  5;
            Y_COORD_14_58_1: value  <=  6;
            Y_COORD_14_59_0: value  <=  9;
            Y_COORD_14_59_1: value  <=  9;
            Y_COORD_14_60_0: value  <=  9;
            Y_COORD_14_60_1: value  <=  9;
            Y_COORD_14_61_0: value  <=  17;
            Y_COORD_14_61_1: value  <=  18;
            Y_COORD_14_62_0: value  <=  16;
            Y_COORD_14_62_1: value  <=  16;
            Y_COORD_14_62_2: value  <=  18;
            Y_COORD_14_63_0: value  <=  16;
            Y_COORD_14_63_1: value  <=  17;
            Y_COORD_14_64_0: value  <=  13;
            Y_COORD_14_64_1: value  <=  15;
            Y_COORD_14_65_0: value  <=  14;
            Y_COORD_14_65_1: value  <=  17;
            Y_COORD_14_66_0: value  <=  15;
            Y_COORD_14_66_1: value  <=  16;
            Y_COORD_14_67_0: value  <=  10;
            Y_COORD_14_67_1: value  <=  12;
            Y_COORD_14_68_0: value  <=  11;
            Y_COORD_14_68_1: value  <=  12;
            Y_COORD_14_69_0: value  <=  9;
            Y_COORD_14_69_1: value  <=  10;
            Y_COORD_14_70_0: value  <=  8;
            Y_COORD_14_70_1: value  <=  9;
            Y_COORD_14_71_0: value  <=  5;
            Y_COORD_14_71_1: value  <=  5;
            Y_COORD_14_72_0: value  <=  19;
            Y_COORD_14_72_1: value  <=  19;
            Y_COORD_14_73_0: value  <=  0;
            Y_COORD_14_73_1: value  <=  0;
            Y_COORD_14_74_0: value  <=  8;
            Y_COORD_14_74_1: value  <=  10;
            Y_COORD_14_75_0: value  <=  17;
            Y_COORD_14_75_1: value  <=  17;
            Y_COORD_14_76_0: value  <=  5;
            Y_COORD_14_76_1: value  <=  5;
            Y_COORD_14_77_0: value  <=  7;
            Y_COORD_14_77_1: value  <=  8;
            Y_COORD_14_78_0: value  <=  11;
            Y_COORD_14_78_1: value  <=  11;
            Y_COORD_14_78_2: value  <=  12;
            Y_COORD_14_79_0: value  <=  3;
            Y_COORD_14_79_1: value  <=  3;
            Y_COORD_14_80_0: value  <=  3;
            Y_COORD_14_80_1: value  <=  3;
            Y_COORD_14_81_0: value  <=  13;
            Y_COORD_14_81_1: value  <=  14;
            Y_COORD_14_82_0: value  <=  6;
            Y_COORD_14_82_1: value  <=  7;
            Y_COORD_14_83_0: value  <=  19;
            Y_COORD_14_83_1: value  <=  19;
            Y_COORD_14_84_0: value  <=  19;
            Y_COORD_14_84_1: value  <=  19;
            Y_COORD_14_85_0: value  <=  13;
            Y_COORD_14_85_1: value  <=  14;
            Y_COORD_14_86_0: value  <=  0;
            Y_COORD_14_86_1: value  <=  0;
            Y_COORD_14_87_0: value  <=  6;
            Y_COORD_14_87_1: value  <=  6;
            Y_COORD_14_88_0: value  <=  5;
            Y_COORD_14_88_1: value  <=  5;
            Y_COORD_14_89_0: value  <=  11;
            Y_COORD_14_89_1: value  <=  12;
            Y_COORD_14_90_0: value  <=  11;
            Y_COORD_14_90_1: value  <=  12;
            Y_COORD_14_91_0: value  <=  6;
            Y_COORD_14_91_1: value  <=  7;
            Y_COORD_14_92_0: value  <=  15;
            Y_COORD_14_92_1: value  <=  16;
            Y_COORD_14_93_0: value  <=  0;
            Y_COORD_14_93_1: value  <=  0;
            Y_COORD_14_94_0: value  <=  0;
            Y_COORD_14_94_1: value  <=  0;
            Y_COORD_14_95_0: value  <=  10;
            Y_COORD_14_95_1: value  <=  10;
            Y_COORD_14_95_2: value  <=  15;
            Y_COORD_14_96_0: value  <=  2;
            Y_COORD_14_96_1: value  <=  2;
            Y_COORD_14_97_0: value  <=  2;
            Y_COORD_14_97_1: value  <=  3;
            Y_COORD_14_98_0: value  <=  10;
            Y_COORD_14_98_1: value  <=  10;
            Y_COORD_14_98_2: value  <=  15;
            Y_COORD_14_99_0: value  <=  13;
            Y_COORD_14_99_1: value  <=  13;
            Y_COORD_14_99_2: value  <=  16;
            Y_COORD_14_100_0: value  <=  5;
            Y_COORD_14_100_1: value  <=  5;
            Y_COORD_14_101_0: value  <=  7;
            Y_COORD_14_101_1: value  <=  7;
            Y_COORD_14_101_2: value  <=  9;
            Y_COORD_14_102_0: value  <=  0;
            Y_COORD_14_102_1: value  <=  0;
            Y_COORD_14_103_0: value  <=  6;
            Y_COORD_14_103_1: value  <=  6;
            Y_COORD_14_103_2: value  <=  9;
            Y_COORD_14_104_0: value  <=  14;
            Y_COORD_14_104_1: value  <=  15;
            Y_COORD_14_105_0: value  <=  15;
            Y_COORD_14_105_1: value  <=  16;
            Y_COORD_14_106_0: value  <=  2;
            Y_COORD_14_106_1: value  <=  2;
            Y_COORD_14_106_2: value  <=  3;
            Y_COORD_14_107_0: value  <=  11;
            Y_COORD_14_107_1: value  <=  14;
            Y_COORD_14_108_0: value  <=  13;
            Y_COORD_14_108_1: value  <=  14;
            Y_COORD_14_109_0: value  <=  4;
            Y_COORD_14_109_1: value  <=  6;
            Y_COORD_14_110_0: value  <=  12;
            Y_COORD_14_110_1: value  <=  13;
            Y_COORD_14_111_0: value  <=  4;
            Y_COORD_14_111_1: value  <=  6;
            Y_COORD_14_112_0: value  <=  13;
            Y_COORD_14_112_1: value  <=  14;
            Y_COORD_14_113_0: value  <=  4;
            Y_COORD_14_113_1: value  <=  6;
            Y_COORD_14_114_0: value  <=  4;
            Y_COORD_14_114_1: value  <=  6;
            Y_COORD_14_115_0: value  <=  12;
            Y_COORD_14_115_1: value  <=  13;
            Y_COORD_14_116_0: value  <=  13;
            Y_COORD_14_116_1: value  <=  14;
            Y_COORD_14_117_0: value  <=  13;
            Y_COORD_14_117_1: value  <=  14;
            Y_COORD_14_118_0: value  <=  4;
            Y_COORD_14_118_1: value  <=  5;
            Y_COORD_14_119_0: value  <=  2;
            Y_COORD_14_119_1: value  <=  4;
            Y_COORD_14_120_0: value  <=  13;
            Y_COORD_14_120_1: value  <=  14;
            Y_COORD_14_121_0: value  <=  7;
            Y_COORD_14_121_1: value  <=  7;
            Y_COORD_14_122_0: value  <=  7;
            Y_COORD_14_122_1: value  <=  7;
            Y_COORD_14_123_0: value  <=  3;
            Y_COORD_14_123_1: value  <=  3;
            Y_COORD_14_124_0: value  <=  6;
            Y_COORD_14_124_1: value  <=  6;
            Y_COORD_14_125_0: value  <=  7;
            Y_COORD_14_125_1: value  <=  8;
            Y_COORD_14_126_0: value  <=  9;
            Y_COORD_14_126_1: value  <=  9;
            Y_COORD_14_127_0: value  <=  13;
            Y_COORD_14_127_1: value  <=  13;
            Y_COORD_14_128_0: value  <=  7;
            Y_COORD_14_128_1: value  <=  7;
            Y_COORD_14_129_0: value  <=  7;
            Y_COORD_14_129_1: value  <=  7;
            Y_COORD_14_130_0: value  <=  7;
            Y_COORD_14_130_1: value  <=  7;
            Y_COORD_14_131_0: value  <=  9;
            Y_COORD_14_131_1: value  <=  9;
            Y_COORD_14_132_0: value  <=  6;
            Y_COORD_14_132_1: value  <=  6;
            Y_COORD_14_133_0: value  <=  12;
            Y_COORD_14_133_1: value  <=  12;
            Y_COORD_14_134_0: value  <=  1;
            Y_COORD_14_134_1: value  <=  6;
            Y_COORD_15_0_0: value  <=  0;
            Y_COORD_15_0_1: value  <=  0;
            Y_COORD_15_1_0: value  <=  7;
            Y_COORD_15_1_1: value  <=  7;
            Y_COORD_15_2_0: value  <=  16;
            Y_COORD_15_2_1: value  <=  16;
            Y_COORD_15_2_2: value  <=  18;
            Y_COORD_15_3_0: value  <=  5;
            Y_COORD_15_3_1: value  <=  9;
            Y_COORD_15_4_0: value  <=  10;
            Y_COORD_15_4_1: value  <=  13;
            Y_COORD_15_5_0: value  <=  6;
            Y_COORD_15_5_1: value  <=  6;
            Y_COORD_15_5_2: value  <=  11;
            Y_COORD_15_6_0: value  <=  6;
            Y_COORD_15_6_1: value  <=  6;
            Y_COORD_15_6_2: value  <=  11;
            Y_COORD_15_7_0: value  <=  5;
            Y_COORD_15_7_1: value  <=  6;
            Y_COORD_15_8_0: value  <=  12;
            Y_COORD_15_8_1: value  <=  13;
            Y_COORD_15_9_0: value  <=  2;
            Y_COORD_15_9_1: value  <=  3;
            Y_COORD_15_10_0: value  <=  0;
            Y_COORD_15_10_1: value  <=  0;
            Y_COORD_15_10_2: value  <=  5;
            Y_COORD_15_11_0: value  <=  10;
            Y_COORD_15_11_1: value  <=  11;
            Y_COORD_15_12_0: value  <=  8;
            Y_COORD_15_12_1: value  <=  9;
            Y_COORD_15_13_0: value  <=  13;
            Y_COORD_15_13_1: value  <=  14;
            Y_COORD_15_14_0: value  <=  2;
            Y_COORD_15_14_1: value  <=  2;
            Y_COORD_15_15_0: value  <=  13;
            Y_COORD_15_15_1: value  <=  14;
            Y_COORD_15_16_0: value  <=  9;
            Y_COORD_15_16_1: value  <=  10;
            Y_COORD_15_17_0: value  <=  2;
            Y_COORD_15_17_1: value  <=  4;
            Y_COORD_15_18_0: value  <=  5;
            Y_COORD_15_18_1: value  <=  5;
            Y_COORD_15_19_0: value  <=  8;
            Y_COORD_15_19_1: value  <=  10;
            Y_COORD_15_20_0: value  <=  4;
            Y_COORD_15_20_1: value  <=  4;
            Y_COORD_15_21_0: value  <=  13;
            Y_COORD_15_21_1: value  <=  16;
            Y_COORD_15_22_0: value  <=  14;
            Y_COORD_15_22_1: value  <=  15;
            Y_COORD_15_23_0: value  <=  8;
            Y_COORD_15_23_1: value  <=  10;
            Y_COORD_15_24_0: value  <=  8;
            Y_COORD_15_24_1: value  <=  10;
            Y_COORD_15_25_0: value  <=  14;
            Y_COORD_15_25_1: value  <=  17;
            Y_COORD_15_26_0: value  <=  5;
            Y_COORD_15_26_1: value  <=  5;
            Y_COORD_15_27_0: value  <=  2;
            Y_COORD_15_27_1: value  <=  2;
            Y_COORD_15_27_2: value  <=  5;
            Y_COORD_15_28_0: value  <=  6;
            Y_COORD_15_28_1: value  <=  6;
            Y_COORD_15_29_0: value  <=  1;
            Y_COORD_15_29_1: value  <=  3;
            Y_COORD_15_30_0: value  <=  7;
            Y_COORD_15_30_1: value  <=  7;
            Y_COORD_15_31_0: value  <=  18;
            Y_COORD_15_31_1: value  <=  18;
            Y_COORD_15_32_0: value  <=  18;
            Y_COORD_15_32_1: value  <=  18;
            Y_COORD_15_33_0: value  <=  3;
            Y_COORD_15_33_1: value  <=  4;
            Y_COORD_15_34_0: value  <=  1;
            Y_COORD_15_34_1: value  <=  7;
            Y_COORD_15_35_0: value  <=  0;
            Y_COORD_15_35_1: value  <=  0;
            Y_COORD_15_36_0: value  <=  2;
            Y_COORD_15_36_1: value  <=  3;
            Y_COORD_15_37_0: value  <=  14;
            Y_COORD_15_37_1: value  <=  14;
            Y_COORD_15_37_2: value  <=  15;
            Y_COORD_15_38_0: value  <=  2;
            Y_COORD_15_38_1: value  <=  4;
            Y_COORD_15_39_0: value  <=  7;
            Y_COORD_15_39_1: value  <=  8;
            Y_COORD_15_40_0: value  <=  5;
            Y_COORD_15_40_1: value  <=  6;
            Y_COORD_15_41_0: value  <=  10;
            Y_COORD_15_41_1: value  <=  10;
            Y_COORD_15_42_0: value  <=  10;
            Y_COORD_15_42_1: value  <=  10;
            Y_COORD_15_43_0: value  <=  17;
            Y_COORD_15_43_1: value  <=  18;
            Y_COORD_15_44_0: value  <=  14;
            Y_COORD_15_44_1: value  <=  15;
            Y_COORD_15_45_0: value  <=  5;
            Y_COORD_15_45_1: value  <=  6;
            Y_COORD_15_46_0: value  <=  5;
            Y_COORD_15_46_1: value  <=  6;
            Y_COORD_15_47_0: value  <=  8;
            Y_COORD_15_47_1: value  <=  9;
            Y_COORD_15_48_0: value  <=  9;
            Y_COORD_15_48_1: value  <=  9;
            Y_COORD_15_49_0: value  <=  0;
            Y_COORD_15_49_1: value  <=  0;
            Y_COORD_15_50_0: value  <=  12;
            Y_COORD_15_50_1: value  <=  13;
            Y_COORD_15_51_0: value  <=  5;
            Y_COORD_15_51_1: value  <=  10;
            Y_COORD_15_52_0: value  <=  14;
            Y_COORD_15_52_1: value  <=  15;
            Y_COORD_15_53_0: value  <=  14;
            Y_COORD_15_53_1: value  <=  15;
            Y_COORD_15_54_0: value  <=  1;
            Y_COORD_15_54_1: value  <=  1;
            Y_COORD_15_55_0: value  <=  0;
            Y_COORD_15_55_1: value  <=  0;
            Y_COORD_15_56_0: value  <=  13;
            Y_COORD_15_56_1: value  <=  14;
            Y_COORD_15_57_0: value  <=  11;
            Y_COORD_15_57_1: value  <=  12;
            Y_COORD_15_58_0: value  <=  5;
            Y_COORD_15_58_1: value  <=  10;
            Y_COORD_15_59_0: value  <=  0;
            Y_COORD_15_59_1: value  <=  0;
            Y_COORD_15_59_2: value  <=  5;
            Y_COORD_15_60_0: value  <=  1;
            Y_COORD_15_60_1: value  <=  1;
            Y_COORD_15_61_0: value  <=  7;
            Y_COORD_15_61_1: value  <=  7;
            Y_COORD_15_62_0: value  <=  1;
            Y_COORD_15_62_1: value  <=  1;
            Y_COORD_15_62_2: value  <=  6;
            Y_COORD_15_63_0: value  <=  7;
            Y_COORD_15_63_1: value  <=  7;
            Y_COORD_15_64_0: value  <=  13;
            Y_COORD_15_64_1: value  <=  15;
            Y_COORD_15_65_0: value  <=  7;
            Y_COORD_15_65_1: value  <=  7;
            Y_COORD_15_66_0: value  <=  7;
            Y_COORD_15_66_1: value  <=  7;
            Y_COORD_15_67_0: value  <=  12;
            Y_COORD_15_67_1: value  <=  12;
            Y_COORD_15_67_2: value  <=  14;
            Y_COORD_15_68_0: value  <=  7;
            Y_COORD_15_68_1: value  <=  7;
            Y_COORD_15_68_2: value  <=  8;
            Y_COORD_15_69_0: value  <=  3;
            Y_COORD_15_69_1: value  <=  4;
            Y_COORD_15_70_0: value  <=  2;
            Y_COORD_15_70_1: value  <=  2;
            Y_COORD_15_70_2: value  <=  11;
            Y_COORD_15_71_0: value  <=  2;
            Y_COORD_15_71_1: value  <=  2;
            Y_COORD_15_71_2: value  <=  4;
            Y_COORD_15_72_0: value  <=  14;
            Y_COORD_15_72_1: value  <=  15;
            Y_COORD_15_73_0: value  <=  12;
            Y_COORD_15_73_1: value  <=  12;
            Y_COORD_15_73_2: value  <=  14;
            Y_COORD_15_74_0: value  <=  12;
            Y_COORD_15_74_1: value  <=  12;
            Y_COORD_15_74_2: value  <=  14;
            Y_COORD_15_75_0: value  <=  4;
            Y_COORD_15_75_1: value  <=  5;
            Y_COORD_15_76_0: value  <=  4;
            Y_COORD_15_76_1: value  <=  5;
            Y_COORD_15_77_0: value  <=  17;
            Y_COORD_15_77_1: value  <=  18;
            Y_COORD_15_78_0: value  <=  1;
            Y_COORD_15_78_1: value  <=  1;
            Y_COORD_15_79_0: value  <=  4;
            Y_COORD_15_79_1: value  <=  4;
            Y_COORD_15_80_0: value  <=  17;
            Y_COORD_15_80_1: value  <=  17;
            Y_COORD_15_81_0: value  <=  0;
            Y_COORD_15_81_1: value  <=  0;
            Y_COORD_15_81_2: value  <=  4;
            Y_COORD_15_82_0: value  <=  8;
            Y_COORD_15_82_1: value  <=  8;
            Y_COORD_15_82_2: value  <=  14;
            Y_COORD_15_83_0: value  <=  7;
            Y_COORD_15_83_1: value  <=  13;
            Y_COORD_15_84_0: value  <=  3;
            Y_COORD_15_84_1: value  <=  10;
            Y_COORD_15_85_0: value  <=  10;
            Y_COORD_15_85_1: value  <=  10;
            Y_COORD_15_86_0: value  <=  4;
            Y_COORD_15_86_1: value  <=  6;
            Y_COORD_15_87_0: value  <=  0;
            Y_COORD_15_87_1: value  <=  4;
            Y_COORD_15_88_0: value  <=  1;
            Y_COORD_15_88_1: value  <=  1;
            Y_COORD_15_88_2: value  <=  5;
            Y_COORD_15_89_0: value  <=  11;
            Y_COORD_15_89_1: value  <=  11;
            Y_COORD_15_90_0: value  <=  9;
            Y_COORD_15_90_1: value  <=  9;
            Y_COORD_15_91_0: value  <=  4;
            Y_COORD_15_91_1: value  <=  6;
            Y_COORD_15_92_0: value  <=  8;
            Y_COORD_15_92_1: value  <=  8;
            Y_COORD_15_93_0: value  <=  1;
            Y_COORD_15_93_1: value  <=  2;
            Y_COORD_15_94_0: value  <=  13;
            Y_COORD_15_94_1: value  <=  13;
            Y_COORD_15_95_0: value  <=  11;
            Y_COORD_15_95_1: value  <=  13;
            Y_COORD_15_96_0: value  <=  11;
            Y_COORD_15_96_1: value  <=  11;
            Y_COORD_15_97_0: value  <=  4;
            Y_COORD_15_97_1: value  <=  4;
            Y_COORD_15_97_2: value  <=  9;
            Y_COORD_15_98_0: value  <=  6;
            Y_COORD_15_98_1: value  <=  9;
            Y_COORD_15_99_0: value  <=  6;
            Y_COORD_15_99_1: value  <=  7;
            Y_COORD_15_100_0: value  <=  7;
            Y_COORD_15_100_1: value  <=  7;
            Y_COORD_15_101_0: value  <=  15;
            Y_COORD_15_101_1: value  <=  16;
            Y_COORD_15_102_0: value  <=  10;
            Y_COORD_15_102_1: value  <=  10;
            Y_COORD_15_103_0: value  <=  15;
            Y_COORD_15_103_1: value  <=  16;
            Y_COORD_15_104_0: value  <=  8;
            Y_COORD_15_104_1: value  <=  10;
            Y_COORD_15_105_0: value  <=  15;
            Y_COORD_15_105_1: value  <=  16;
            Y_COORD_15_106_0: value  <=  15;
            Y_COORD_15_106_1: value  <=  16;
            Y_COORD_15_107_0: value  <=  3;
            Y_COORD_15_107_1: value  <=  3;
            Y_COORD_15_107_2: value  <=  7;
            Y_COORD_15_108_0: value  <=  3;
            Y_COORD_15_108_1: value  <=  3;
            Y_COORD_15_108_2: value  <=  7;
            Y_COORD_15_109_0: value  <=  7;
            Y_COORD_15_109_1: value  <=  7;
            Y_COORD_15_109_2: value  <=  12;
            Y_COORD_15_110_0: value  <=  7;
            Y_COORD_15_110_1: value  <=  8;
            Y_COORD_15_111_0: value  <=  6;
            Y_COORD_15_111_1: value  <=  7;
            Y_COORD_15_112_0: value  <=  6;
            Y_COORD_15_112_1: value  <=  7;
            Y_COORD_15_113_0: value  <=  6;
            Y_COORD_15_113_1: value  <=  7;
            Y_COORD_15_114_0: value  <=  6;
            Y_COORD_15_114_1: value  <=  7;
            Y_COORD_15_115_0: value  <=  2;
            Y_COORD_15_115_1: value  <=  3;
            Y_COORD_15_116_0: value  <=  3;
            Y_COORD_15_116_1: value  <=  3;
            Y_COORD_15_117_0: value  <=  6;
            Y_COORD_15_117_1: value  <=  7;
            Y_COORD_15_118_0: value  <=  10;
            Y_COORD_15_118_1: value  <=  12;
            Y_COORD_15_119_0: value  <=  0;
            Y_COORD_15_119_1: value  <=  7;
            Y_COORD_15_120_0: value  <=  0;
            Y_COORD_15_120_1: value  <=  0;
            Y_COORD_15_120_2: value  <=  5;
            Y_COORD_15_121_0: value  <=  6;
            Y_COORD_15_121_1: value  <=  6;
            Y_COORD_15_122_0: value  <=  6;
            Y_COORD_15_122_1: value  <=  6;
            Y_COORD_15_123_0: value  <=  2;
            Y_COORD_15_123_1: value  <=  3;
            Y_COORD_15_124_0: value  <=  2;
            Y_COORD_15_124_1: value  <=  3;
            Y_COORD_15_125_0: value  <=  11;
            Y_COORD_15_125_1: value  <=  11;
            Y_COORD_15_125_2: value  <=  12;
            Y_COORD_15_126_0: value  <=  5;
            Y_COORD_15_126_1: value  <=  5;
            Y_COORD_15_126_2: value  <=  6;
            Y_COORD_15_127_0: value  <=  9;
            Y_COORD_15_127_1: value  <=  9;
            Y_COORD_15_128_0: value  <=  1;
            Y_COORD_15_128_1: value  <=  1;
            Y_COORD_15_129_0: value  <=  4;
            Y_COORD_15_129_1: value  <=  5;
            Y_COORD_15_130_0: value  <=  4;
            Y_COORD_15_130_1: value  <=  5;
            Y_COORD_15_131_0: value  <=  5;
            Y_COORD_15_131_1: value  <=  6;
            Y_COORD_15_132_0: value  <=  16;
            Y_COORD_15_132_1: value  <=  17;
            Y_COORD_15_133_0: value  <=  13;
            Y_COORD_15_133_1: value  <=  13;
            Y_COORD_15_133_2: value  <=  16;
            Y_COORD_15_134_0: value  <=  5;
            Y_COORD_15_134_1: value  <=  6;
            Y_COORD_15_135_0: value  <=  0;
            Y_COORD_15_135_1: value  <=  0;
            Y_COORD_15_136_0: value  <=  1;
            Y_COORD_15_136_1: value  <=  1;
            Y_COORD_15_136_2: value  <=  4;
            Y_COORD_16_0_0: value  <=  4;
            Y_COORD_16_0_1: value  <=  6;
            Y_COORD_16_1_0: value  <=  2;
            Y_COORD_16_1_1: value  <=  2;
            Y_COORD_16_2_0: value  <=  6;
            Y_COORD_16_2_1: value  <=  12;
            Y_COORD_16_3_0: value  <=  5;
            Y_COORD_16_3_1: value  <=  9;
            Y_COORD_16_4_0: value  <=  4;
            Y_COORD_16_4_1: value  <=  4;
            Y_COORD_16_4_2: value  <=  9;
            Y_COORD_16_5_0: value  <=  6;
            Y_COORD_16_5_1: value  <=  6;
            Y_COORD_16_5_2: value  <=  13;
            Y_COORD_16_6_0: value  <=  6;
            Y_COORD_16_6_1: value  <=  6;
            Y_COORD_16_6_2: value  <=  13;
            Y_COORD_16_7_0: value  <=  9;
            Y_COORD_16_7_1: value  <=  9;
            Y_COORD_16_8_0: value  <=  14;
            Y_COORD_16_8_1: value  <=  15;
            Y_COORD_16_9_0: value  <=  3;
            Y_COORD_16_9_1: value  <=  3;
            Y_COORD_16_9_2: value  <=  5;
            Y_COORD_16_10_0: value  <=  9;
            Y_COORD_16_10_1: value  <=  9;
            Y_COORD_16_11_0: value  <=  11;
            Y_COORD_16_11_1: value  <=  14;
            Y_COORD_16_12_0: value  <=  4;
            Y_COORD_16_12_1: value  <=  4;
            Y_COORD_16_13_0: value  <=  6;
            Y_COORD_16_13_1: value  <=  9;
            Y_COORD_16_14_0: value  <=  7;
            Y_COORD_16_14_1: value  <=  7;
            Y_COORD_16_14_2: value  <=  9;
            Y_COORD_16_15_0: value  <=  1;
            Y_COORD_16_15_1: value  <=  1;
            Y_COORD_16_16_0: value  <=  2;
            Y_COORD_16_16_1: value  <=  2;
            Y_COORD_16_17_0: value  <=  17;
            Y_COORD_16_17_1: value  <=  18;
            Y_COORD_16_18_0: value  <=  17;
            Y_COORD_16_18_1: value  <=  18;
            Y_COORD_16_19_0: value  <=  3;
            Y_COORD_16_19_1: value  <=  5;
            Y_COORD_16_20_0: value  <=  17;
            Y_COORD_16_20_1: value  <=  18;
            Y_COORD_16_21_0: value  <=  13;
            Y_COORD_16_21_1: value  <=  16;
            Y_COORD_16_22_0: value  <=  13;
            Y_COORD_16_22_1: value  <=  14;
            Y_COORD_16_23_0: value  <=  3;
            Y_COORD_16_23_1: value  <=  5;
            Y_COORD_16_24_0: value  <=  13;
            Y_COORD_16_24_1: value  <=  14;
            Y_COORD_16_25_0: value  <=  3;
            Y_COORD_16_25_1: value  <=  3;
            Y_COORD_16_26_0: value  <=  3;
            Y_COORD_16_26_1: value  <=  5;
            Y_COORD_16_27_0: value  <=  5;
            Y_COORD_16_27_1: value  <=  7;
            Y_COORD_16_28_0: value  <=  5;
            Y_COORD_16_28_1: value  <=  6;
            Y_COORD_16_29_0: value  <=  1;
            Y_COORD_16_29_1: value  <=  1;
            Y_COORD_16_30_0: value  <=  2;
            Y_COORD_16_30_1: value  <=  5;
            Y_COORD_16_31_0: value  <=  6;
            Y_COORD_16_31_1: value  <=  7;
            Y_COORD_16_32_0: value  <=  6;
            Y_COORD_16_32_1: value  <=  6;
            Y_COORD_16_33_0: value  <=  11;
            Y_COORD_16_33_1: value  <=  15;
            Y_COORD_16_34_0: value  <=  6;
            Y_COORD_16_34_1: value  <=  7;
            Y_COORD_16_35_0: value  <=  6;
            Y_COORD_16_35_1: value  <=  6;
            Y_COORD_16_35_2: value  <=  7;
            Y_COORD_16_36_0: value  <=  6;
            Y_COORD_16_36_1: value  <=  6;
            Y_COORD_16_36_2: value  <=  7;
            Y_COORD_16_37_0: value  <=  1;
            Y_COORD_16_37_1: value  <=  1;
            Y_COORD_16_38_0: value  <=  1;
            Y_COORD_16_38_1: value  <=  1;
            Y_COORD_16_39_0: value  <=  2;
            Y_COORD_16_39_1: value  <=  9;
            Y_COORD_16_40_0: value  <=  7;
            Y_COORD_16_40_1: value  <=  7;
            Y_COORD_16_41_0: value  <=  3;
            Y_COORD_16_41_1: value  <=  3;
            Y_COORD_16_41_2: value  <=  5;
            Y_COORD_16_42_0: value  <=  7;
            Y_COORD_16_42_1: value  <=  7;
            Y_COORD_16_43_0: value  <=  9;
            Y_COORD_16_43_1: value  <=  9;
            Y_COORD_16_44_0: value  <=  2;
            Y_COORD_16_44_1: value  <=  2;
            Y_COORD_16_45_0: value  <=  5;
            Y_COORD_16_45_1: value  <=  5;
            Y_COORD_16_46_0: value  <=  9;
            Y_COORD_16_46_1: value  <=  9;
            Y_COORD_16_47_0: value  <=  0;
            Y_COORD_16_47_1: value  <=  9;
            Y_COORD_16_48_0: value  <=  16;
            Y_COORD_16_48_1: value  <=  17;
            Y_COORD_16_49_0: value  <=  7;
            Y_COORD_16_49_1: value  <=  7;
            Y_COORD_16_50_0: value  <=  8;
            Y_COORD_16_50_1: value  <=  9;
            Y_COORD_16_51_0: value  <=  12;
            Y_COORD_16_51_1: value  <=  13;
            Y_COORD_16_52_0: value  <=  12;
            Y_COORD_16_52_1: value  <=  13;
            Y_COORD_16_53_0: value  <=  12;
            Y_COORD_16_53_1: value  <=  12;
            Y_COORD_16_54_0: value  <=  11;
            Y_COORD_16_54_1: value  <=  14;
            Y_COORD_16_55_0: value  <=  12;
            Y_COORD_16_55_1: value  <=  13;
            Y_COORD_16_56_0: value  <=  10;
            Y_COORD_16_56_1: value  <=  10;
            Y_COORD_16_56_2: value  <=  13;
            Y_COORD_16_57_0: value  <=  10;
            Y_COORD_16_57_1: value  <=  12;
            Y_COORD_16_58_0: value  <=  16;
            Y_COORD_16_58_1: value  <=  17;
            Y_COORD_16_59_0: value  <=  3;
            Y_COORD_16_59_1: value  <=  6;
            Y_COORD_16_60_0: value  <=  13;
            Y_COORD_16_60_1: value  <=  15;
            Y_COORD_16_61_0: value  <=  6;
            Y_COORD_16_61_1: value  <=  9;
            Y_COORD_16_62_0: value  <=  4;
            Y_COORD_16_62_1: value  <=  4;
            Y_COORD_16_63_0: value  <=  0;
            Y_COORD_16_63_1: value  <=  0;
            Y_COORD_16_64_0: value  <=  3;
            Y_COORD_16_64_1: value  <=  4;
            Y_COORD_16_65_0: value  <=  0;
            Y_COORD_16_65_1: value  <=  2;
            Y_COORD_16_66_0: value  <=  6;
            Y_COORD_16_66_1: value  <=  9;
            Y_COORD_16_67_0: value  <=  8;
            Y_COORD_16_67_1: value  <=  9;
            Y_COORD_16_68_0: value  <=  0;
            Y_COORD_16_68_1: value  <=  0;
            Y_COORD_16_69_0: value  <=  18;
            Y_COORD_16_69_1: value  <=  18;
            Y_COORD_16_69_2: value  <=  19;
            Y_COORD_16_70_0: value  <=  15;
            Y_COORD_16_70_1: value  <=  16;
            Y_COORD_16_71_0: value  <=  14;
            Y_COORD_16_71_1: value  <=  15;
            Y_COORD_16_72_0: value  <=  14;
            Y_COORD_16_72_1: value  <=  15;
            Y_COORD_16_73_0: value  <=  3;
            Y_COORD_16_73_1: value  <=  3;
            Y_COORD_16_74_0: value  <=  5;
            Y_COORD_16_74_1: value  <=  5;
            Y_COORD_16_75_0: value  <=  5;
            Y_COORD_16_75_1: value  <=  6;
            Y_COORD_16_76_0: value  <=  5;
            Y_COORD_16_76_1: value  <=  6;
            Y_COORD_16_77_0: value  <=  14;
            Y_COORD_16_77_1: value  <=  17;
            Y_COORD_16_78_0: value  <=  9;
            Y_COORD_16_78_1: value  <=  9;
            Y_COORD_16_79_0: value  <=  3;
            Y_COORD_16_79_1: value  <=  3;
            Y_COORD_16_80_0: value  <=  0;
            Y_COORD_16_80_1: value  <=  0;
            Y_COORD_16_81_0: value  <=  6;
            Y_COORD_16_81_1: value  <=  7;
            Y_COORD_16_82_0: value  <=  14;
            Y_COORD_16_82_1: value  <=  17;
            Y_COORD_16_83_0: value  <=  8;
            Y_COORD_16_83_1: value  <=  9;
            Y_COORD_16_84_0: value  <=  3;
            Y_COORD_16_84_1: value  <=  3;
            Y_COORD_16_85_0: value  <=  16;
            Y_COORD_16_85_1: value  <=  17;
            Y_COORD_16_86_0: value  <=  6;
            Y_COORD_16_86_1: value  <=  7;
            Y_COORD_16_87_0: value  <=  4;
            Y_COORD_16_87_1: value  <=  4;
            Y_COORD_16_87_2: value  <=  5;
            Y_COORD_16_88_0: value  <=  4;
            Y_COORD_16_88_1: value  <=  4;
            Y_COORD_16_88_2: value  <=  5;
            Y_COORD_16_89_0: value  <=  16;
            Y_COORD_16_89_1: value  <=  18;
            Y_COORD_16_90_0: value  <=  15;
            Y_COORD_16_90_1: value  <=  17;
            Y_COORD_16_91_0: value  <=  0;
            Y_COORD_16_91_1: value  <=  1;
            Y_COORD_16_92_0: value  <=  0;
            Y_COORD_16_92_1: value  <=  0;
            Y_COORD_16_93_0: value  <=  4;
            Y_COORD_16_93_1: value  <=  4;
            Y_COORD_16_93_2: value  <=  8;
            Y_COORD_16_94_0: value  <=  7;
            Y_COORD_16_94_1: value  <=  7;
            Y_COORD_16_94_2: value  <=  8;
            Y_COORD_16_95_0: value  <=  6;
            Y_COORD_16_95_1: value  <=  7;
            Y_COORD_16_96_0: value  <=  7;
            Y_COORD_16_96_1: value  <=  8;
            Y_COORD_16_97_0: value  <=  2;
            Y_COORD_16_97_1: value  <=  8;
            Y_COORD_16_98_0: value  <=  0;
            Y_COORD_16_98_1: value  <=  4;
            Y_COORD_16_99_0: value  <=  9;
            Y_COORD_16_99_1: value  <=  9;
            Y_COORD_16_100_0: value  <=  14;
            Y_COORD_16_100_1: value  <=  15;
            Y_COORD_16_101_0: value  <=  10;
            Y_COORD_16_101_1: value  <=  11;
            Y_COORD_16_102_0: value  <=  11;
            Y_COORD_16_102_1: value  <=  12;
            Y_COORD_16_103_0: value  <=  15;
            Y_COORD_16_103_1: value  <=  15;
            Y_COORD_16_104_0: value  <=  8;
            Y_COORD_16_104_1: value  <=  8;
            Y_COORD_16_105_0: value  <=  15;
            Y_COORD_16_105_1: value  <=  15;
            Y_COORD_16_106_0: value  <=  7;
            Y_COORD_16_106_1: value  <=  7;
            Y_COORD_16_107_0: value  <=  10;
            Y_COORD_16_107_1: value  <=  10;
            Y_COORD_16_107_2: value  <=  12;
            Y_COORD_16_108_0: value  <=  3;
            Y_COORD_16_108_1: value  <=  3;
            Y_COORD_16_109_0: value  <=  13;
            Y_COORD_16_109_1: value  <=  13;
            Y_COORD_16_110_0: value  <=  2;
            Y_COORD_16_110_1: value  <=  2;
            Y_COORD_16_111_0: value  <=  2;
            Y_COORD_16_111_1: value  <=  2;
            Y_COORD_16_112_0: value  <=  0;
            Y_COORD_16_112_1: value  <=  0;
            Y_COORD_16_112_2: value  <=  6;
            Y_COORD_16_113_0: value  <=  7;
            Y_COORD_16_113_1: value  <=  7;
            Y_COORD_16_113_2: value  <=  8;
            Y_COORD_16_114_0: value  <=  12;
            Y_COORD_16_114_1: value  <=  14;
            Y_COORD_16_115_0: value  <=  7;
            Y_COORD_16_115_1: value  <=  7;
            Y_COORD_16_116_0: value  <=  8;
            Y_COORD_16_116_1: value  <=  8;
            Y_COORD_16_117_0: value  <=  0;
            Y_COORD_16_117_1: value  <=  0;
            Y_COORD_16_118_0: value  <=  15;
            Y_COORD_16_118_1: value  <=  16;
            Y_COORD_16_119_0: value  <=  15;
            Y_COORD_16_119_1: value  <=  16;
            Y_COORD_16_120_0: value  <=  10;
            Y_COORD_16_120_1: value  <=  12;
            Y_COORD_16_121_0: value  <=  9;
            Y_COORD_16_121_1: value  <=  10;
            Y_COORD_16_122_0: value  <=  15;
            Y_COORD_16_122_1: value  <=  16;
            Y_COORD_16_123_0: value  <=  7;
            Y_COORD_16_123_1: value  <=  7;
            Y_COORD_16_124_0: value  <=  0;
            Y_COORD_16_124_1: value  <=  0;
            Y_COORD_16_125_0: value  <=  6;
            Y_COORD_16_125_1: value  <=  6;
            Y_COORD_16_125_2: value  <=  9;
            Y_COORD_16_126_0: value  <=  6;
            Y_COORD_16_126_1: value  <=  6;
            Y_COORD_16_126_2: value  <=  7;
            Y_COORD_16_127_0: value  <=  6;
            Y_COORD_16_127_1: value  <=  6;
            Y_COORD_16_127_2: value  <=  7;
            Y_COORD_16_128_0: value  <=  6;
            Y_COORD_16_128_1: value  <=  6;
            Y_COORD_16_128_2: value  <=  7;
            Y_COORD_16_129_0: value  <=  4;
            Y_COORD_16_129_1: value  <=  10;
            Y_COORD_16_130_0: value  <=  5;
            Y_COORD_16_130_1: value  <=  5;
            Y_COORD_16_130_2: value  <=  10;
            Y_COORD_16_131_0: value  <=  17;
            Y_COORD_16_131_1: value  <=  17;
            Y_COORD_16_132_0: value  <=  4;
            Y_COORD_16_132_1: value  <=  5;
            Y_COORD_16_133_0: value  <=  0;
            Y_COORD_16_133_1: value  <=  0;
            Y_COORD_16_134_0: value  <=  0;
            Y_COORD_16_134_1: value  <=  0;
            Y_COORD_16_135_0: value  <=  2;
            Y_COORD_16_135_1: value  <=  2;
            Y_COORD_16_136_0: value  <=  2;
            Y_COORD_16_136_1: value  <=  2;
            Y_COORD_16_137_0: value  <=  11;
            Y_COORD_16_137_1: value  <=  11;
            Y_COORD_16_138_0: value  <=  11;
            Y_COORD_16_138_1: value  <=  11;
            Y_COORD_16_139_0: value  <=  16;
            Y_COORD_16_139_1: value  <=  16;
            Y_COORD_17_0_0: value  <=  4;
            Y_COORD_17_0_1: value  <=  4;
            Y_COORD_17_1_0: value  <=  7;
            Y_COORD_17_1_1: value  <=  7;
            Y_COORD_17_1_2: value  <=  9;
            Y_COORD_17_2_0: value  <=  8;
            Y_COORD_17_2_1: value  <=  12;
            Y_COORD_17_3_0: value  <=  1;
            Y_COORD_17_3_1: value  <=  3;
            Y_COORD_17_4_0: value  <=  2;
            Y_COORD_17_4_1: value  <=  2;
            Y_COORD_17_4_2: value  <=  5;
            Y_COORD_17_5_0: value  <=  16;
            Y_COORD_17_5_1: value  <=  16;
            Y_COORD_17_5_2: value  <=  18;
            Y_COORD_17_6_0: value  <=  2;
            Y_COORD_17_6_1: value  <=  2;
            Y_COORD_17_7_0: value  <=  4;
            Y_COORD_17_7_1: value  <=  9;
            Y_COORD_17_8_0: value  <=  9;
            Y_COORD_17_8_1: value  <=  9;
            Y_COORD_17_9_0: value  <=  10;
            Y_COORD_17_9_1: value  <=  13;
            Y_COORD_17_10_0: value  <=  11;
            Y_COORD_17_10_1: value  <=  12;
            Y_COORD_17_11_0: value  <=  11;
            Y_COORD_17_11_1: value  <=  11;
            Y_COORD_17_11_2: value  <=  14;
            Y_COORD_17_12_0: value  <=  0;
            Y_COORD_17_12_1: value  <=  3;
            Y_COORD_17_13_0: value  <=  14;
            Y_COORD_17_13_1: value  <=  16;
            Y_COORD_17_14_0: value  <=  2;
            Y_COORD_17_14_1: value  <=  4;
            Y_COORD_17_15_0: value  <=  14;
            Y_COORD_17_15_1: value  <=  15;
            Y_COORD_17_16_0: value  <=  14;
            Y_COORD_17_16_1: value  <=  16;
            Y_COORD_17_17_0: value  <=  15;
            Y_COORD_17_17_1: value  <=  16;
            Y_COORD_17_18_0: value  <=  4;
            Y_COORD_17_18_1: value  <=  4;
            Y_COORD_17_19_0: value  <=  0;
            Y_COORD_17_19_1: value  <=  1;
            Y_COORD_17_20_0: value  <=  6;
            Y_COORD_17_20_1: value  <=  7;
            Y_COORD_17_21_0: value  <=  1;
            Y_COORD_17_21_1: value  <=  2;
            Y_COORD_17_22_0: value  <=  6;
            Y_COORD_17_22_1: value  <=  6;
            Y_COORD_17_23_0: value  <=  8;
            Y_COORD_17_23_1: value  <=  8;
            Y_COORD_17_24_0: value  <=  8;
            Y_COORD_17_24_1: value  <=  8;
            Y_COORD_17_25_0: value  <=  7;
            Y_COORD_17_25_1: value  <=  7;
            Y_COORD_17_26_0: value  <=  9;
            Y_COORD_17_26_1: value  <=  9;
            Y_COORD_17_27_0: value  <=  9;
            Y_COORD_17_27_1: value  <=  10;
            Y_COORD_17_28_0: value  <=  0;
            Y_COORD_17_28_1: value  <=  0;
            Y_COORD_17_29_0: value  <=  9;
            Y_COORD_17_29_1: value  <=  10;
            Y_COORD_17_30_0: value  <=  10;
            Y_COORD_17_30_1: value  <=  10;
            Y_COORD_17_31_0: value  <=  4;
            Y_COORD_17_31_1: value  <=  4;
            Y_COORD_17_32_0: value  <=  8;
            Y_COORD_17_32_1: value  <=  9;
            Y_COORD_17_33_0: value  <=  2;
            Y_COORD_17_33_1: value  <=  2;
            Y_COORD_17_34_0: value  <=  17;
            Y_COORD_17_34_1: value  <=  18;
            Y_COORD_17_35_0: value  <=  10;
            Y_COORD_17_35_1: value  <=  15;
            Y_COORD_17_36_0: value  <=  7;
            Y_COORD_17_36_1: value  <=  7;
            Y_COORD_17_37_0: value  <=  4;
            Y_COORD_17_37_1: value  <=  4;
            Y_COORD_17_38_0: value  <=  4;
            Y_COORD_17_38_1: value  <=  4;
            Y_COORD_17_39_0: value  <=  6;
            Y_COORD_17_39_1: value  <=  6;
            Y_COORD_17_40_0: value  <=  0;
            Y_COORD_17_40_1: value  <=  0;
            Y_COORD_17_40_2: value  <=  6;
            Y_COORD_17_41_0: value  <=  2;
            Y_COORD_17_41_1: value  <=  2;
            Y_COORD_17_42_0: value  <=  0;
            Y_COORD_17_42_1: value  <=  0;
            Y_COORD_17_43_0: value  <=  2;
            Y_COORD_17_43_1: value  <=  2;
            Y_COORD_17_44_0: value  <=  5;
            Y_COORD_17_44_1: value  <=  8;
            Y_COORD_17_45_0: value  <=  12;
            Y_COORD_17_45_1: value  <=  12;
            Y_COORD_17_45_2: value  <=  13;
            Y_COORD_17_46_0: value  <=  17;
            Y_COORD_17_46_1: value  <=  17;
            Y_COORD_17_47_0: value  <=  6;
            Y_COORD_17_47_1: value  <=  6;
            Y_COORD_17_47_2: value  <=  7;
            Y_COORD_17_48_0: value  <=  9;
            Y_COORD_17_48_1: value  <=  9;
            Y_COORD_17_49_0: value  <=  6;
            Y_COORD_17_49_1: value  <=  6;
            Y_COORD_17_49_2: value  <=  7;
            Y_COORD_17_50_0: value  <=  4;
            Y_COORD_17_50_1: value  <=  4;
            Y_COORD_17_51_0: value  <=  11;
            Y_COORD_17_51_1: value  <=  12;
            Y_COORD_17_52_0: value  <=  10;
            Y_COORD_17_52_1: value  <=  11;
            Y_COORD_17_53_0: value  <=  7;
            Y_COORD_17_53_1: value  <=  7;
            Y_COORD_17_54_0: value  <=  4;
            Y_COORD_17_54_1: value  <=  5;
            Y_COORD_17_55_0: value  <=  4;
            Y_COORD_17_55_1: value  <=  5;
            Y_COORD_17_56_0: value  <=  4;
            Y_COORD_17_56_1: value  <=  5;
            Y_COORD_17_57_0: value  <=  8;
            Y_COORD_17_57_1: value  <=  9;
            Y_COORD_17_58_0: value  <=  9;
            Y_COORD_17_58_1: value  <=  10;
            Y_COORD_17_59_0: value  <=  14;
            Y_COORD_17_59_1: value  <=  16;
            Y_COORD_17_60_0: value  <=  12;
            Y_COORD_17_60_1: value  <=  13;
            Y_COORD_17_61_0: value  <=  15;
            Y_COORD_17_61_1: value  <=  15;
            Y_COORD_17_61_2: value  <=  16;
            Y_COORD_17_62_0: value  <=  13;
            Y_COORD_17_62_1: value  <=  14;
            Y_COORD_17_63_0: value  <=  11;
            Y_COORD_17_63_1: value  <=  14;
            Y_COORD_17_64_0: value  <=  13;
            Y_COORD_17_64_1: value  <=  14;
            Y_COORD_17_65_0: value  <=  14;
            Y_COORD_17_65_1: value  <=  16;
            Y_COORD_17_66_0: value  <=  14;
            Y_COORD_17_66_1: value  <=  16;
            Y_COORD_17_67_0: value  <=  0;
            Y_COORD_17_67_1: value  <=  0;
            Y_COORD_17_68_0: value  <=  1;
            Y_COORD_17_68_1: value  <=  1;
            Y_COORD_17_68_2: value  <=  7;
            Y_COORD_17_69_0: value  <=  14;
            Y_COORD_17_69_1: value  <=  14;
            Y_COORD_17_69_2: value  <=  17;
            Y_COORD_17_70_0: value  <=  14;
            Y_COORD_17_70_1: value  <=  14;
            Y_COORD_17_70_2: value  <=  17;
            Y_COORD_17_71_0: value  <=  17;
            Y_COORD_17_71_1: value  <=  18;
            Y_COORD_17_72_0: value  <=  17;
            Y_COORD_17_72_1: value  <=  18;
            Y_COORD_17_73_0: value  <=  0;
            Y_COORD_17_73_1: value  <=  0;
            Y_COORD_17_74_0: value  <=  0;
            Y_COORD_17_74_1: value  <=  0;
            Y_COORD_17_75_0: value  <=  10;
            Y_COORD_17_75_1: value  <=  12;
            Y_COORD_17_76_0: value  <=  15;
            Y_COORD_17_76_1: value  <=  15;
            Y_COORD_17_76_2: value  <=  16;
            Y_COORD_17_77_0: value  <=  11;
            Y_COORD_17_77_1: value  <=  11;
            Y_COORD_17_77_2: value  <=  14;
            Y_COORD_17_78_0: value  <=  6;
            Y_COORD_17_78_1: value  <=  6;
            Y_COORD_17_78_2: value  <=  7;
            Y_COORD_17_79_0: value  <=  2;
            Y_COORD_17_79_1: value  <=  2;
            Y_COORD_17_79_2: value  <=  5;
            Y_COORD_17_80_0: value  <=  4;
            Y_COORD_17_80_1: value  <=  5;
            Y_COORD_17_81_0: value  <=  7;
            Y_COORD_17_81_1: value  <=  12;
            Y_COORD_17_82_0: value  <=  7;
            Y_COORD_17_82_1: value  <=  12;
            Y_COORD_17_83_0: value  <=  7;
            Y_COORD_17_83_1: value  <=  7;
            Y_COORD_17_84_0: value  <=  12;
            Y_COORD_17_84_1: value  <=  13;
            Y_COORD_17_85_0: value  <=  1;
            Y_COORD_17_85_1: value  <=  2;
            Y_COORD_17_86_0: value  <=  2;
            Y_COORD_17_86_1: value  <=  2;
            Y_COORD_17_86_2: value  <=  11;
            Y_COORD_17_87_0: value  <=  4;
            Y_COORD_17_87_1: value  <=  10;
            Y_COORD_17_88_0: value  <=  0;
            Y_COORD_17_88_1: value  <=  2;
            Y_COORD_17_89_0: value  <=  11;
            Y_COORD_17_89_1: value  <=  12;
            Y_COORD_17_90_0: value  <=  7;
            Y_COORD_17_90_1: value  <=  8;
            Y_COORD_17_91_0: value  <=  7;
            Y_COORD_17_91_1: value  <=  7;
            Y_COORD_17_92_0: value  <=  7;
            Y_COORD_17_92_1: value  <=  7;
            Y_COORD_17_93_0: value  <=  4;
            Y_COORD_17_93_1: value  <=  4;
            Y_COORD_17_94_0: value  <=  7;
            Y_COORD_17_94_1: value  <=  7;
            Y_COORD_17_95_0: value  <=  7;
            Y_COORD_17_95_1: value  <=  7;
            Y_COORD_17_95_2: value  <=  10;
            Y_COORD_17_96_0: value  <=  7;
            Y_COORD_17_96_1: value  <=  7;
            Y_COORD_17_96_2: value  <=  10;
            Y_COORD_17_97_0: value  <=  2;
            Y_COORD_17_97_1: value  <=  2;
            Y_COORD_17_97_2: value  <=  7;
            Y_COORD_17_98_0: value  <=  2;
            Y_COORD_17_98_1: value  <=  2;
            Y_COORD_17_99_0: value  <=  4;
            Y_COORD_17_99_1: value  <=  4;
            Y_COORD_17_100_0: value  <=  15;
            Y_COORD_17_100_1: value  <=  15;
            Y_COORD_17_100_2: value  <=  16;
            Y_COORD_17_101_0: value  <=  13;
            Y_COORD_17_101_1: value  <=  16;
            Y_COORD_17_102_0: value  <=  13;
            Y_COORD_17_102_1: value  <=  16;
            Y_COORD_17_103_0: value  <=  3;
            Y_COORD_17_103_1: value  <=  3;
            Y_COORD_17_104_0: value  <=  15;
            Y_COORD_17_104_1: value  <=  16;
            Y_COORD_17_105_0: value  <=  15;
            Y_COORD_17_105_1: value  <=  17;
            Y_COORD_17_106_0: value  <=  14;
            Y_COORD_17_106_1: value  <=  15;
            Y_COORD_17_107_0: value  <=  3;
            Y_COORD_17_107_1: value  <=  3;
            Y_COORD_17_108_0: value  <=  12;
            Y_COORD_17_108_1: value  <=  13;
            Y_COORD_17_109_0: value  <=  11;
            Y_COORD_17_109_1: value  <=  14;
            Y_COORD_17_110_0: value  <=  13;
            Y_COORD_17_110_1: value  <=  13;
            Y_COORD_17_110_2: value  <=  14;
            Y_COORD_17_111_0: value  <=  11;
            Y_COORD_17_111_1: value  <=  11;
            Y_COORD_17_111_2: value  <=  13;
            Y_COORD_17_112_0: value  <=  18;
            Y_COORD_17_112_1: value  <=  18;
            Y_COORD_17_113_0: value  <=  18;
            Y_COORD_17_113_1: value  <=  18;
            Y_COORD_17_113_2: value  <=  19;
            Y_COORD_17_114_0: value  <=  18;
            Y_COORD_17_114_1: value  <=  18;
            Y_COORD_17_114_2: value  <=  19;
            Y_COORD_17_115_0: value  <=  18;
            Y_COORD_17_115_1: value  <=  19;
            Y_COORD_17_116_0: value  <=  14;
            Y_COORD_17_116_1: value  <=  15;
            Y_COORD_17_117_0: value  <=  12;
            Y_COORD_17_117_1: value  <=  12;
            Y_COORD_17_117_2: value  <=  16;
            Y_COORD_17_118_0: value  <=  9;
            Y_COORD_17_118_1: value  <=  10;
            Y_COORD_17_119_0: value  <=  10;
            Y_COORD_17_119_1: value  <=  10;
            Y_COORD_17_120_0: value  <=  0;
            Y_COORD_17_120_1: value  <=  0;
            Y_COORD_17_121_0: value  <=  6;
            Y_COORD_17_121_1: value  <=  6;
            Y_COORD_17_122_0: value  <=  16;
            Y_COORD_17_122_1: value  <=  17;
            Y_COORD_17_123_0: value  <=  1;
            Y_COORD_17_123_1: value  <=  1;
            Y_COORD_17_124_0: value  <=  0;
            Y_COORD_17_124_1: value  <=  1;
            Y_COORD_17_125_0: value  <=  12;
            Y_COORD_17_125_1: value  <=  12;
            Y_COORD_17_126_0: value  <=  12;
            Y_COORD_17_126_1: value  <=  12;
            Y_COORD_17_127_0: value  <=  11;
            Y_COORD_17_127_1: value  <=  11;
            Y_COORD_17_127_2: value  <=  12;
            Y_COORD_17_128_0: value  <=  2;
            Y_COORD_17_128_1: value  <=  4;
            Y_COORD_17_129_0: value  <=  11;
            Y_COORD_17_129_1: value  <=  11;
            Y_COORD_17_129_2: value  <=  12;
            Y_COORD_17_130_0: value  <=  6;
            Y_COORD_17_130_1: value  <=  11;
            Y_COORD_17_131_0: value  <=  11;
            Y_COORD_17_131_1: value  <=  11;
            Y_COORD_17_131_2: value  <=  12;
            Y_COORD_17_132_0: value  <=  13;
            Y_COORD_17_132_1: value  <=  14;
            Y_COORD_17_133_0: value  <=  11;
            Y_COORD_17_133_1: value  <=  11;
            Y_COORD_17_133_2: value  <=  12;
            Y_COORD_17_134_0: value  <=  11;
            Y_COORD_17_134_1: value  <=  11;
            Y_COORD_17_134_2: value  <=  12;
            Y_COORD_17_135_0: value  <=  13;
            Y_COORD_17_135_1: value  <=  14;
            Y_COORD_17_136_0: value  <=  13;
            Y_COORD_17_136_1: value  <=  14;
            Y_COORD_17_137_0: value  <=  14;
            Y_COORD_17_137_1: value  <=  15;
            Y_COORD_17_138_0: value  <=  7;
            Y_COORD_17_138_1: value  <=  8;
            Y_COORD_17_139_0: value  <=  5;
            Y_COORD_17_139_1: value  <=  6;
            Y_COORD_17_140_0: value  <=  9;
            Y_COORD_17_140_1: value  <=  10;
            Y_COORD_17_141_0: value  <=  5;
            Y_COORD_17_141_1: value  <=  6;
            Y_COORD_17_142_0: value  <=  12;
            Y_COORD_17_142_1: value  <=  12;
            Y_COORD_17_142_2: value  <=  16;
            Y_COORD_17_143_0: value  <=  7;
            Y_COORD_17_143_1: value  <=  7;
            Y_COORD_17_143_2: value  <=  8;
            Y_COORD_17_144_0: value  <=  16;
            Y_COORD_17_144_1: value  <=  16;
            Y_COORD_17_145_0: value  <=  6;
            Y_COORD_17_145_1: value  <=  7;
            Y_COORD_17_146_0: value  <=  5;
            Y_COORD_17_146_1: value  <=  7;
            Y_COORD_17_147_0: value  <=  15;
            Y_COORD_17_147_1: value  <=  15;
            Y_COORD_17_148_0: value  <=  14;
            Y_COORD_17_148_1: value  <=  14;
            Y_COORD_17_149_0: value  <=  0;
            Y_COORD_17_149_1: value  <=  0;
            Y_COORD_17_150_0: value  <=  15;
            Y_COORD_17_150_1: value  <=  15;
            Y_COORD_17_151_0: value  <=  7;
            Y_COORD_17_151_1: value  <=  7;
            Y_COORD_17_152_0: value  <=  7;
            Y_COORD_17_152_1: value  <=  7;
            Y_COORD_17_153_0: value  <=  6;
            Y_COORD_17_153_1: value  <=  9;
            Y_COORD_17_154_0: value  <=  4;
            Y_COORD_17_154_1: value  <=  10;
            Y_COORD_17_155_0: value  <=  12;
            Y_COORD_17_155_1: value  <=  12;
            Y_COORD_17_155_2: value  <=  13;
            Y_COORD_17_156_0: value  <=  12;
            Y_COORD_17_156_1: value  <=  12;
            Y_COORD_17_156_2: value  <=  13;
            Y_COORD_17_157_0: value  <=  9;
            Y_COORD_17_157_1: value  <=  9;
            Y_COORD_17_157_2: value  <=  10;
            Y_COORD_17_158_0: value  <=  6;
            Y_COORD_17_158_1: value  <=  6;
            Y_COORD_17_158_2: value  <=  7;
            Y_COORD_17_159_0: value  <=  6;
            Y_COORD_17_159_1: value  <=  7;
            Y_COORD_18_0_0: value  <=  7;
            Y_COORD_18_0_1: value  <=  9;
            Y_COORD_18_1_0: value  <=  2;
            Y_COORD_18_1_1: value  <=  2;
            Y_COORD_18_2_0: value  <=  4;
            Y_COORD_18_2_1: value  <=  10;
            Y_COORD_18_3_0: value  <=  18;
            Y_COORD_18_3_1: value  <=  18;
            Y_COORD_18_4_0: value  <=  7;
            Y_COORD_18_4_1: value  <=  7;
            Y_COORD_18_4_2: value  <=  9;
            Y_COORD_18_5_0: value  <=  0;
            Y_COORD_18_5_1: value  <=  0;
            Y_COORD_18_6_0: value  <=  0;
            Y_COORD_18_6_1: value  <=  0;
            Y_COORD_18_7_0: value  <=  5;
            Y_COORD_18_7_1: value  <=  9;
            Y_COORD_18_8_0: value  <=  3;
            Y_COORD_18_8_1: value  <=  3;
            Y_COORD_18_9_0: value  <=  4;
            Y_COORD_18_9_1: value  <=  4;
            Y_COORD_18_10_0: value  <=  4;
            Y_COORD_18_10_1: value  <=  4;
            Y_COORD_18_11_0: value  <=  0;
            Y_COORD_18_11_1: value  <=  0;
            Y_COORD_18_12_0: value  <=  17;
            Y_COORD_18_12_1: value  <=  18;
            Y_COORD_18_13_0: value  <=  11;
            Y_COORD_18_13_1: value  <=  11;
            Y_COORD_18_14_0: value  <=  2;
            Y_COORD_18_14_1: value  <=  3;
            Y_COORD_18_15_0: value  <=  12;
            Y_COORD_18_15_1: value  <=  13;
            Y_COORD_18_16_0: value  <=  10;
            Y_COORD_18_16_1: value  <=  13;
            Y_COORD_18_17_0: value  <=  4;
            Y_COORD_18_17_1: value  <=  4;
            Y_COORD_18_18_0: value  <=  4;
            Y_COORD_18_18_1: value  <=  4;
            Y_COORD_18_19_0: value  <=  6;
            Y_COORD_18_19_1: value  <=  6;
            Y_COORD_18_20_0: value  <=  13;
            Y_COORD_18_20_1: value  <=  14;
            Y_COORD_18_21_0: value  <=  15;
            Y_COORD_18_21_1: value  <=  15;
            Y_COORD_18_22_0: value  <=  2;
            Y_COORD_18_22_1: value  <=  2;
            Y_COORD_18_23_0: value  <=  0;
            Y_COORD_18_23_1: value  <=  0;
            Y_COORD_18_24_0: value  <=  15;
            Y_COORD_18_24_1: value  <=  15;
            Y_COORD_18_25_0: value  <=  13;
            Y_COORD_18_25_1: value  <=  14;
            Y_COORD_18_26_0: value  <=  16;
            Y_COORD_18_26_1: value  <=  16;
            Y_COORD_18_27_0: value  <=  2;
            Y_COORD_18_27_1: value  <=  7;
            Y_COORD_18_28_0: value  <=  5;
            Y_COORD_18_28_1: value  <=  9;
            Y_COORD_18_29_0: value  <=  16;
            Y_COORD_18_29_1: value  <=  17;
            Y_COORD_18_30_0: value  <=  16;
            Y_COORD_18_30_1: value  <=  17;
            Y_COORD_18_31_0: value  <=  11;
            Y_COORD_18_31_1: value  <=  14;
            Y_COORD_18_32_0: value  <=  11;
            Y_COORD_18_32_1: value  <=  14;
            Y_COORD_18_33_0: value  <=  14;
            Y_COORD_18_33_1: value  <=  15;
            Y_COORD_18_34_0: value  <=  14;
            Y_COORD_18_34_1: value  <=  15;
            Y_COORD_18_35_0: value  <=  0;
            Y_COORD_18_35_1: value  <=  0;
            Y_COORD_18_35_2: value  <=  3;
            Y_COORD_18_36_0: value  <=  3;
            Y_COORD_18_36_1: value  <=  4;
            Y_COORD_18_37_0: value  <=  0;
            Y_COORD_18_37_1: value  <=  0;
            Y_COORD_18_37_2: value  <=  1;
            Y_COORD_18_38_0: value  <=  12;
            Y_COORD_18_38_1: value  <=  16;
            Y_COORD_18_39_0: value  <=  7;
            Y_COORD_18_39_1: value  <=  7;
            Y_COORD_18_39_2: value  <=  12;
            Y_COORD_18_40_0: value  <=  7;
            Y_COORD_18_40_1: value  <=  7;
            Y_COORD_18_40_2: value  <=  12;
            Y_COORD_18_41_0: value  <=  10;
            Y_COORD_18_41_1: value  <=  12;
            Y_COORD_18_42_0: value  <=  4;
            Y_COORD_18_42_1: value  <=  4;
            Y_COORD_18_43_0: value  <=  5;
            Y_COORD_18_43_1: value  <=  7;
            Y_COORD_18_44_0: value  <=  0;
            Y_COORD_18_44_1: value  <=  0;
            Y_COORD_18_44_2: value  <=  1;
            Y_COORD_18_45_0: value  <=  0;
            Y_COORD_18_45_1: value  <=  0;
            Y_COORD_18_46_0: value  <=  13;
            Y_COORD_18_46_1: value  <=  14;
            Y_COORD_18_47_0: value  <=  8;
            Y_COORD_18_47_1: value  <=  8;
            Y_COORD_18_48_0: value  <=  1;
            Y_COORD_18_48_1: value  <=  1;
            Y_COORD_18_49_0: value  <=  14;
            Y_COORD_18_49_1: value  <=  15;
            Y_COORD_18_50_0: value  <=  6;
            Y_COORD_18_50_1: value  <=  6;
            Y_COORD_18_51_0: value  <=  11;
            Y_COORD_18_51_1: value  <=  12;
            Y_COORD_18_52_0: value  <=  5;
            Y_COORD_18_52_1: value  <=  6;
            Y_COORD_18_53_0: value  <=  4;
            Y_COORD_18_53_1: value  <=  5;
            Y_COORD_18_54_0: value  <=  15;
            Y_COORD_18_54_1: value  <=  16;
            Y_COORD_18_55_0: value  <=  4;
            Y_COORD_18_55_1: value  <=  5;
            Y_COORD_18_56_0: value  <=  0;
            Y_COORD_18_56_1: value  <=  1;
            Y_COORD_18_57_0: value  <=  12;
            Y_COORD_18_57_1: value  <=  12;
            Y_COORD_18_58_0: value  <=  4;
            Y_COORD_18_58_1: value  <=  5;
            Y_COORD_18_59_0: value  <=  4;
            Y_COORD_18_59_1: value  <=  5;
            Y_COORD_18_60_0: value  <=  0;
            Y_COORD_18_60_1: value  <=  2;
            Y_COORD_18_61_0: value  <=  2;
            Y_COORD_18_61_1: value  <=  2;
            Y_COORD_18_61_2: value  <=  5;
            Y_COORD_18_62_0: value  <=  7;
            Y_COORD_18_62_1: value  <=  7;
            Y_COORD_18_63_0: value  <=  10;
            Y_COORD_18_63_1: value  <=  10;
            Y_COORD_18_64_0: value  <=  0;
            Y_COORD_18_64_1: value  <=  0;
            Y_COORD_18_65_0: value  <=  0;
            Y_COORD_18_65_1: value  <=  0;
            Y_COORD_18_66_0: value  <=  19;
            Y_COORD_18_66_1: value  <=  19;
            Y_COORD_18_67_0: value  <=  10;
            Y_COORD_18_67_1: value  <=  10;
            Y_COORD_18_67_2: value  <=  15;
            Y_COORD_18_68_0: value  <=  8;
            Y_COORD_18_68_1: value  <=  9;
            Y_COORD_18_69_0: value  <=  12;
            Y_COORD_18_69_1: value  <=  13;
            Y_COORD_18_70_0: value  <=  10;
            Y_COORD_18_70_1: value  <=  10;
            Y_COORD_18_70_2: value  <=  15;
            Y_COORD_18_71_0: value  <=  3;
            Y_COORD_18_71_1: value  <=  5;
            Y_COORD_18_72_0: value  <=  6;
            Y_COORD_18_72_1: value  <=  7;
            Y_COORD_18_73_0: value  <=  7;
            Y_COORD_18_73_1: value  <=  8;
            Y_COORD_18_74_0: value  <=  3;
            Y_COORD_18_74_1: value  <=  5;
            Y_COORD_18_75_0: value  <=  1;
            Y_COORD_18_75_1: value  <=  1;
            Y_COORD_18_76_0: value  <=  0;
            Y_COORD_18_76_1: value  <=  0;
            Y_COORD_18_77_0: value  <=  1;
            Y_COORD_18_77_1: value  <=  1;
            Y_COORD_18_78_0: value  <=  6;
            Y_COORD_18_78_1: value  <=  6;
            Y_COORD_18_79_0: value  <=  12;
            Y_COORD_18_79_1: value  <=  12;
            Y_COORD_18_80_0: value  <=  12;
            Y_COORD_18_80_1: value  <=  12;
            Y_COORD_18_81_0: value  <=  7;
            Y_COORD_18_81_1: value  <=  7;
            Y_COORD_18_82_0: value  <=  7;
            Y_COORD_18_82_1: value  <=  7;
            Y_COORD_18_83_0: value  <=  0;
            Y_COORD_18_83_1: value  <=  0;
            Y_COORD_18_84_0: value  <=  11;
            Y_COORD_18_84_1: value  <=  12;
            Y_COORD_18_85_0: value  <=  3;
            Y_COORD_18_85_1: value  <=  3;
            Y_COORD_18_86_0: value  <=  8;
            Y_COORD_18_86_1: value  <=  13;
            Y_COORD_18_87_0: value  <=  0;
            Y_COORD_18_87_1: value  <=  0;
            Y_COORD_18_88_0: value  <=  14;
            Y_COORD_18_88_1: value  <=  15;
            Y_COORD_18_89_0: value  <=  3;
            Y_COORD_18_89_1: value  <=  3;
            Y_COORD_18_90_0: value  <=  0;
            Y_COORD_18_90_1: value  <=  0;
            Y_COORD_18_91_0: value  <=  3;
            Y_COORD_18_91_1: value  <=  3;
            Y_COORD_18_92_0: value  <=  9;
            Y_COORD_18_92_1: value  <=  10;
            Y_COORD_18_93_0: value  <=  1;
            Y_COORD_18_93_1: value  <=  1;
            Y_COORD_18_94_0: value  <=  1;
            Y_COORD_18_94_1: value  <=  1;
            Y_COORD_18_95_0: value  <=  16;
            Y_COORD_18_95_1: value  <=  16;
            Y_COORD_18_96_0: value  <=  8;
            Y_COORD_18_96_1: value  <=  8;
            Y_COORD_18_97_0: value  <=  0;
            Y_COORD_18_97_1: value  <=  0;
            Y_COORD_18_97_2: value  <=  3;
            Y_COORD_18_98_0: value  <=  0;
            Y_COORD_18_98_1: value  <=  0;
            Y_COORD_18_98_2: value  <=  3;
            Y_COORD_18_99_0: value  <=  3;
            Y_COORD_18_99_1: value  <=  3;
            Y_COORD_18_100_0: value  <=  3;
            Y_COORD_18_100_1: value  <=  3;
            Y_COORD_18_101_0: value  <=  1;
            Y_COORD_18_101_1: value  <=  1;
            Y_COORD_18_102_0: value  <=  1;
            Y_COORD_18_102_1: value  <=  1;
            Y_COORD_18_103_0: value  <=  0;
            Y_COORD_18_103_1: value  <=  0;
            Y_COORD_18_103_2: value  <=  4;
            Y_COORD_18_104_0: value  <=  8;
            Y_COORD_18_104_1: value  <=  9;
            Y_COORD_18_105_0: value  <=  7;
            Y_COORD_18_105_1: value  <=  7;
            Y_COORD_18_106_0: value  <=  8;
            Y_COORD_18_106_1: value  <=  9;
            Y_COORD_18_107_0: value  <=  6;
            Y_COORD_18_107_1: value  <=  6;
            Y_COORD_18_108_0: value  <=  7;
            Y_COORD_18_108_1: value  <=  7;
            Y_COORD_18_109_0: value  <=  2;
            Y_COORD_18_109_1: value  <=  5;
            Y_COORD_18_110_0: value  <=  7;
            Y_COORD_18_110_1: value  <=  7;
            Y_COORD_18_110_2: value  <=  9;
            Y_COORD_18_111_0: value  <=  12;
            Y_COORD_18_111_1: value  <=  13;
            Y_COORD_18_112_0: value  <=  11;
            Y_COORD_18_112_1: value  <=  12;
            Y_COORD_18_113_0: value  <=  5;
            Y_COORD_18_113_1: value  <=  5;
            Y_COORD_18_113_2: value  <=  10;
            Y_COORD_18_114_0: value  <=  12;
            Y_COORD_18_114_1: value  <=  13;
            Y_COORD_18_115_0: value  <=  11;
            Y_COORD_18_115_1: value  <=  11;
            Y_COORD_18_116_0: value  <=  9;
            Y_COORD_18_116_1: value  <=  11;
            Y_COORD_18_117_0: value  <=  10;
            Y_COORD_18_117_1: value  <=  11;
            Y_COORD_18_118_0: value  <=  11;
            Y_COORD_18_118_1: value  <=  12;
            Y_COORD_18_119_0: value  <=  5;
            Y_COORD_18_119_1: value  <=  7;
            Y_COORD_18_120_0: value  <=  4;
            Y_COORD_18_120_1: value  <=  4;
            Y_COORD_18_121_0: value  <=  11;
            Y_COORD_18_121_1: value  <=  11;
            Y_COORD_18_122_0: value  <=  11;
            Y_COORD_18_122_1: value  <=  11;
            Y_COORD_18_123_0: value  <=  16;
            Y_COORD_18_123_1: value  <=  16;
            Y_COORD_18_124_0: value  <=  7;
            Y_COORD_18_124_1: value  <=  7;
            Y_COORD_18_125_0: value  <=  12;
            Y_COORD_18_125_1: value  <=  16;
            Y_COORD_18_126_0: value  <=  15;
            Y_COORD_18_126_1: value  <=  16;
            Y_COORD_18_127_0: value  <=  4;
            Y_COORD_18_127_1: value  <=  6;
            Y_COORD_18_128_0: value  <=  5;
            Y_COORD_18_128_1: value  <=  5;
            Y_COORD_18_129_0: value  <=  10;
            Y_COORD_18_129_1: value  <=  12;
            Y_COORD_18_130_0: value  <=  19;
            Y_COORD_18_130_1: value  <=  19;
            Y_COORD_18_131_0: value  <=  16;
            Y_COORD_18_131_1: value  <=  16;
            Y_COORD_18_132_0: value  <=  15;
            Y_COORD_18_132_1: value  <=  17;
            Y_COORD_18_133_0: value  <=  16;
            Y_COORD_18_133_1: value  <=  16;
            Y_COORD_18_134_0: value  <=  16;
            Y_COORD_18_134_1: value  <=  16;
            Y_COORD_18_135_0: value  <=  16;
            Y_COORD_18_135_1: value  <=  17;
            Y_COORD_18_136_0: value  <=  11;
            Y_COORD_18_136_1: value  <=  14;
            Y_COORD_18_137_0: value  <=  6;
            Y_COORD_18_137_1: value  <=  10;
            Y_COORD_18_138_0: value  <=  17;
            Y_COORD_18_138_1: value  <=  18;
            Y_COORD_18_139_0: value  <=  18;
            Y_COORD_18_139_1: value  <=  18;
            Y_COORD_18_139_2: value  <=  19;
            Y_COORD_18_140_0: value  <=  18;
            Y_COORD_18_140_1: value  <=  19;
            Y_COORD_18_141_0: value  <=  5;
            Y_COORD_18_141_1: value  <=  5;
            Y_COORD_18_142_0: value  <=  8;
            Y_COORD_18_142_1: value  <=  9;
            Y_COORD_18_143_0: value  <=  5;
            Y_COORD_18_143_1: value  <=  5;
            Y_COORD_18_144_0: value  <=  5;
            Y_COORD_18_144_1: value  <=  5;
            Y_COORD_18_145_0: value  <=  1;
            Y_COORD_18_145_1: value  <=  1;
            Y_COORD_18_145_2: value  <=  5;
            Y_COORD_18_146_0: value  <=  4;
            Y_COORD_18_146_1: value  <=  4;
            Y_COORD_18_146_2: value  <=  12;
            Y_COORD_18_147_0: value  <=  4;
            Y_COORD_18_147_1: value  <=  10;
            Y_COORD_18_148_0: value  <=  5;
            Y_COORD_18_148_1: value  <=  5;
            Y_COORD_18_148_2: value  <=  11;
            Y_COORD_18_149_0: value  <=  14;
            Y_COORD_18_149_1: value  <=  15;
            Y_COORD_18_150_0: value  <=  4;
            Y_COORD_18_150_1: value  <=  5;
            Y_COORD_18_151_0: value  <=  2;
            Y_COORD_18_151_1: value  <=  2;
            Y_COORD_18_151_2: value  <=  7;
            Y_COORD_18_152_0: value  <=  4;
            Y_COORD_18_152_1: value  <=  5;
            Y_COORD_18_153_0: value  <=  0;
            Y_COORD_18_153_1: value  <=  0;
            Y_COORD_18_153_2: value  <=  1;
            Y_COORD_18_154_0: value  <=  0;
            Y_COORD_18_154_1: value  <=  0;
            Y_COORD_18_154_2: value  <=  1;
            Y_COORD_18_155_0: value  <=  13;
            Y_COORD_18_155_1: value  <=  13;
            Y_COORD_18_155_2: value  <=  16;
            Y_COORD_18_156_0: value  <=  13;
            Y_COORD_18_156_1: value  <=  13;
            Y_COORD_18_156_2: value  <=  16;
            Y_COORD_18_157_0: value  <=  12;
            Y_COORD_18_157_1: value  <=  15;
            Y_COORD_18_158_0: value  <=  9;
            Y_COORD_18_158_1: value  <=  9;
            Y_COORD_18_158_2: value  <=  14;
            Y_COORD_18_159_0: value  <=  4;
            Y_COORD_18_159_1: value  <=  4;
            Y_COORD_18_159_2: value  <=  5;
            Y_COORD_18_160_0: value  <=  12;
            Y_COORD_18_160_1: value  <=  12;
            Y_COORD_18_161_0: value  <=  2;
            Y_COORD_18_161_1: value  <=  2;
            Y_COORD_18_161_2: value  <=  7;
            Y_COORD_18_162_0: value  <=  11;
            Y_COORD_18_162_1: value  <=  11;
            Y_COORD_18_163_0: value  <=  5;
            Y_COORD_18_163_1: value  <=  9;
            Y_COORD_18_164_0: value  <=  11;
            Y_COORD_18_164_1: value  <=  11;
            Y_COORD_18_165_0: value  <=  2;
            Y_COORD_18_165_1: value  <=  2;
            Y_COORD_18_165_2: value  <=  7;
            Y_COORD_18_166_0: value  <=  2;
            Y_COORD_18_166_1: value  <=  2;
            Y_COORD_18_166_2: value  <=  7;
            Y_COORD_18_167_0: value  <=  4;
            Y_COORD_18_167_1: value  <=  4;
            Y_COORD_18_167_2: value  <=  5;
            Y_COORD_18_168_0: value  <=  14;
            Y_COORD_18_168_1: value  <=  15;
            Y_COORD_18_169_0: value  <=  4;
            Y_COORD_18_169_1: value  <=  4;
            Y_COORD_18_169_2: value  <=  5;
            Y_COORD_18_170_0: value  <=  1;
            Y_COORD_18_170_1: value  <=  1;
            Y_COORD_18_171_0: value  <=  4;
            Y_COORD_18_171_1: value  <=  4;
            Y_COORD_18_171_2: value  <=  5;
            Y_COORD_18_172_0: value  <=  4;
            Y_COORD_18_172_1: value  <=  4;
            Y_COORD_18_172_2: value  <=  5;
            Y_COORD_18_173_0: value  <=  0;
            Y_COORD_18_173_1: value  <=  0;
            Y_COORD_18_173_2: value  <=  6;
            Y_COORD_18_174_0: value  <=  0;
            Y_COORD_18_174_1: value  <=  0;
            Y_COORD_18_175_0: value  <=  0;
            Y_COORD_18_175_1: value  <=  4;
            Y_COORD_18_176_0: value  <=  4;
            Y_COORD_18_176_1: value  <=  6;
            Y_COORD_19_0_0: value  <=  3;
            Y_COORD_19_0_1: value  <=  3;
            Y_COORD_19_1_0: value  <=  11;
            Y_COORD_19_1_1: value  <=  12;
            Y_COORD_19_2_0: value  <=  7;
            Y_COORD_19_2_1: value  <=  7;
            Y_COORD_19_2_2: value  <=  9;
            Y_COORD_19_3_0: value  <=  3;
            Y_COORD_19_3_1: value  <=  6;
            Y_COORD_19_4_0: value  <=  15;
            Y_COORD_19_4_1: value  <=  17;
            Y_COORD_19_5_0: value  <=  5;
            Y_COORD_19_5_1: value  <=  5;
            Y_COORD_19_6_0: value  <=  2;
            Y_COORD_19_6_1: value  <=  2;
            Y_COORD_19_6_2: value  <=  7;
            Y_COORD_19_7_0: value  <=  0;
            Y_COORD_19_7_1: value  <=  1;
            Y_COORD_19_8_0: value  <=  2;
            Y_COORD_19_8_1: value  <=  7;
            Y_COORD_19_9_0: value  <=  2;
            Y_COORD_19_9_1: value  <=  3;
            Y_COORD_19_10_0: value  <=  3;
            Y_COORD_19_10_1: value  <=  3;
            Y_COORD_19_11_0: value  <=  5;
            Y_COORD_19_11_1: value  <=  10;
            Y_COORD_19_12_0: value  <=  13;
            Y_COORD_19_12_1: value  <=  16;
            Y_COORD_19_13_0: value  <=  7;
            Y_COORD_19_13_1: value  <=  7;
            Y_COORD_19_14_0: value  <=  3;
            Y_COORD_19_14_1: value  <=  3;
            Y_COORD_19_15_0: value  <=  16;
            Y_COORD_19_15_1: value  <=  17;
            Y_COORD_19_16_0: value  <=  2;
            Y_COORD_19_16_1: value  <=  3;
            Y_COORD_19_17_0: value  <=  5;
            Y_COORD_19_17_1: value  <=  6;
            Y_COORD_19_18_0: value  <=  7;
            Y_COORD_19_18_1: value  <=  7;
            Y_COORD_19_19_0: value  <=  5;
            Y_COORD_19_19_1: value  <=  12;
            Y_COORD_19_20_0: value  <=  0;
            Y_COORD_19_20_1: value  <=  0;
            Y_COORD_19_20_2: value  <=  5;
            Y_COORD_19_21_0: value  <=  1;
            Y_COORD_19_21_1: value  <=  1;
            Y_COORD_19_22_0: value  <=  1;
            Y_COORD_19_22_1: value  <=  1;
            Y_COORD_19_23_0: value  <=  4;
            Y_COORD_19_23_1: value  <=  5;
            Y_COORD_19_24_0: value  <=  4;
            Y_COORD_19_24_1: value  <=  12;
            Y_COORD_19_25_0: value  <=  4;
            Y_COORD_19_25_1: value  <=  5;
            Y_COORD_19_26_0: value  <=  3;
            Y_COORD_19_26_1: value  <=  5;
            Y_COORD_19_27_0: value  <=  2;
            Y_COORD_19_27_1: value  <=  5;
            Y_COORD_19_28_0: value  <=  4;
            Y_COORD_19_28_1: value  <=  5;
            Y_COORD_19_29_0: value  <=  17;
            Y_COORD_19_29_1: value  <=  17;
            Y_COORD_19_30_0: value  <=  5;
            Y_COORD_19_30_1: value  <=  6;
            Y_COORD_19_31_0: value  <=  11;
            Y_COORD_19_31_1: value  <=  13;
            Y_COORD_19_32_0: value  <=  14;
            Y_COORD_19_32_1: value  <=  17;
            Y_COORD_19_33_0: value  <=  3;
            Y_COORD_19_33_1: value  <=  4;
            Y_COORD_19_34_0: value  <=  8;
            Y_COORD_19_34_1: value  <=  9;
            Y_COORD_19_35_0: value  <=  3;
            Y_COORD_19_35_1: value  <=  4;
            Y_COORD_19_36_0: value  <=  0;
            Y_COORD_19_36_1: value  <=  2;
            Y_COORD_19_37_0: value  <=  5;
            Y_COORD_19_37_1: value  <=  6;
            Y_COORD_19_38_0: value  <=  11;
            Y_COORD_19_38_1: value  <=  13;
            Y_COORD_19_39_0: value  <=  5;
            Y_COORD_19_39_1: value  <=  6;
            Y_COORD_19_40_0: value  <=  5;
            Y_COORD_19_40_1: value  <=  6;
            Y_COORD_19_41_0: value  <=  5;
            Y_COORD_19_41_1: value  <=  6;
            Y_COORD_19_42_0: value  <=  6;
            Y_COORD_19_42_1: value  <=  12;
            Y_COORD_19_43_0: value  <=  5;
            Y_COORD_19_43_1: value  <=  6;
            Y_COORD_19_44_0: value  <=  12;
            Y_COORD_19_44_1: value  <=  12;
            Y_COORD_19_45_0: value  <=  5;
            Y_COORD_19_45_1: value  <=  6;
            Y_COORD_19_46_0: value  <=  5;
            Y_COORD_19_46_1: value  <=  6;
            Y_COORD_19_47_0: value  <=  6;
            Y_COORD_19_47_1: value  <=  6;
            Y_COORD_19_48_0: value  <=  11;
            Y_COORD_19_48_1: value  <=  12;
            Y_COORD_19_49_0: value  <=  12;
            Y_COORD_19_49_1: value  <=  12;
            Y_COORD_19_50_0: value  <=  0;
            Y_COORD_19_50_1: value  <=  0;
            Y_COORD_19_51_0: value  <=  8;
            Y_COORD_19_51_1: value  <=  8;
            Y_COORD_19_52_0: value  <=  8;
            Y_COORD_19_52_1: value  <=  8;
            Y_COORD_19_53_0: value  <=  10;
            Y_COORD_19_53_1: value  <=  11;
            Y_COORD_19_54_0: value  <=  7;
            Y_COORD_19_54_1: value  <=  7;
            Y_COORD_19_55_0: value  <=  7;
            Y_COORD_19_55_1: value  <=  7;
            Y_COORD_19_56_0: value  <=  7;
            Y_COORD_19_56_1: value  <=  7;
            Y_COORD_19_57_0: value  <=  9;
            Y_COORD_19_57_1: value  <=  9;
            Y_COORD_19_58_0: value  <=  9;
            Y_COORD_19_58_1: value  <=  9;
            Y_COORD_19_59_0: value  <=  10;
            Y_COORD_19_59_1: value  <=  12;
            Y_COORD_19_60_0: value  <=  7;
            Y_COORD_19_60_1: value  <=  7;
            Y_COORD_19_61_0: value  <=  17;
            Y_COORD_19_61_1: value  <=  18;
            Y_COORD_19_62_0: value  <=  5;
            Y_COORD_19_62_1: value  <=  5;
            Y_COORD_19_62_2: value  <=  11;
            Y_COORD_19_63_0: value  <=  9;
            Y_COORD_19_63_1: value  <=  9;
            Y_COORD_19_63_2: value  <=  13;
            Y_COORD_19_64_0: value  <=  4;
            Y_COORD_19_64_1: value  <=  4;
            Y_COORD_19_65_0: value  <=  2;
            Y_COORD_19_65_1: value  <=  2;
            Y_COORD_19_66_0: value  <=  12;
            Y_COORD_19_66_1: value  <=  13;
            Y_COORD_19_67_0: value  <=  13;
            Y_COORD_19_67_1: value  <=  14;
            Y_COORD_19_68_0: value  <=  13;
            Y_COORD_19_68_1: value  <=  14;
            Y_COORD_19_69_0: value  <=  11;
            Y_COORD_19_69_1: value  <=  12;
            Y_COORD_19_70_0: value  <=  12;
            Y_COORD_19_70_1: value  <=  12;
            Y_COORD_19_70_2: value  <=  14;
            Y_COORD_19_71_0: value  <=  11;
            Y_COORD_19_71_1: value  <=  11;
            Y_COORD_19_71_2: value  <=  12;
            Y_COORD_19_72_0: value  <=  17;
            Y_COORD_19_72_1: value  <=  17;
            Y_COORD_19_73_0: value  <=  11;
            Y_COORD_19_73_1: value  <=  11;
            Y_COORD_19_73_2: value  <=  12;
            Y_COORD_19_74_0: value  <=  17;
            Y_COORD_19_74_1: value  <=  18;
            Y_COORD_19_75_0: value  <=  11;
            Y_COORD_19_75_1: value  <=  11;
            Y_COORD_19_75_2: value  <=  12;
            Y_COORD_19_76_0: value  <=  11;
            Y_COORD_19_76_1: value  <=  11;
            Y_COORD_19_76_2: value  <=  12;
            Y_COORD_19_77_0: value  <=  5;
            Y_COORD_19_77_1: value  <=  5;
            Y_COORD_19_78_0: value  <=  5;
            Y_COORD_19_78_1: value  <=  5;
            Y_COORD_19_79_0: value  <=  2;
            Y_COORD_19_79_1: value  <=  2;
            Y_COORD_19_80_0: value  <=  2;
            Y_COORD_19_80_1: value  <=  2;
            Y_COORD_19_81_0: value  <=  0;
            Y_COORD_19_81_1: value  <=  0;
            Y_COORD_19_81_2: value  <=  1;
            Y_COORD_19_82_0: value  <=  12;
            Y_COORD_19_82_1: value  <=  12;
            Y_COORD_19_83_0: value  <=  11;
            Y_COORD_19_83_1: value  <=  11;
            Y_COORD_19_83_2: value  <=  15;
            Y_COORD_19_84_0: value  <=  9;
            Y_COORD_19_84_1: value  <=  10;
            Y_COORD_19_85_0: value  <=  18;
            Y_COORD_19_85_1: value  <=  19;
            Y_COORD_19_86_0: value  <=  6;
            Y_COORD_19_86_1: value  <=  6;
            Y_COORD_19_86_2: value  <=  12;
            Y_COORD_19_87_0: value  <=  8;
            Y_COORD_19_87_1: value  <=  9;
            Y_COORD_19_88_0: value  <=  10;
            Y_COORD_19_88_1: value  <=  10;
            Y_COORD_19_89_0: value  <=  11;
            Y_COORD_19_89_1: value  <=  11;
            Y_COORD_19_90_0: value  <=  11;
            Y_COORD_19_90_1: value  <=  11;
            Y_COORD_19_91_0: value  <=  2;
            Y_COORD_19_91_1: value  <=  2;
            Y_COORD_19_91_2: value  <=  3;
            Y_COORD_19_92_0: value  <=  12;
            Y_COORD_19_92_1: value  <=  13;
            Y_COORD_19_93_0: value  <=  1;
            Y_COORD_19_93_1: value  <=  1;
            Y_COORD_19_94_0: value  <=  1;
            Y_COORD_19_94_1: value  <=  1;
            Y_COORD_19_95_0: value  <=  16;
            Y_COORD_19_95_1: value  <=  16;
            Y_COORD_19_96_0: value  <=  17;
            Y_COORD_19_96_1: value  <=  17;
            Y_COORD_19_97_0: value  <=  14;
            Y_COORD_19_97_1: value  <=  17;
            Y_COORD_19_98_0: value  <=  12;
            Y_COORD_19_98_1: value  <=  16;
            Y_COORD_19_99_0: value  <=  14;
            Y_COORD_19_99_1: value  <=  15;
            Y_COORD_19_100_0: value  <=  6;
            Y_COORD_19_100_1: value  <=  10;
            Y_COORD_19_101_0: value  <=  9;
            Y_COORD_19_101_1: value  <=  10;
            Y_COORD_19_102_0: value  <=  1;
            Y_COORD_19_102_1: value  <=  1;
            Y_COORD_19_103_0: value  <=  1;
            Y_COORD_19_103_1: value  <=  1;
            Y_COORD_19_103_2: value  <=  2;
            Y_COORD_19_104_0: value  <=  3;
            Y_COORD_19_104_1: value  <=  10;
            Y_COORD_19_105_0: value  <=  12;
            Y_COORD_19_105_1: value  <=  12;
            Y_COORD_19_105_2: value  <=  13;
            Y_COORD_19_106_0: value  <=  9;
            Y_COORD_19_106_1: value  <=  9;
            Y_COORD_19_106_2: value  <=  10;
            Y_COORD_19_107_0: value  <=  15;
            Y_COORD_19_107_1: value  <=  16;
            Y_COORD_19_108_0: value  <=  8;
            Y_COORD_19_108_1: value  <=  9;
            Y_COORD_19_109_0: value  <=  15;
            Y_COORD_19_109_1: value  <=  16;
            Y_COORD_19_110_0: value  <=  7;
            Y_COORD_19_110_1: value  <=  8;
            Y_COORD_19_111_0: value  <=  7;
            Y_COORD_19_111_1: value  <=  8;
            Y_COORD_19_112_0: value  <=  7;
            Y_COORD_19_112_1: value  <=  7;
            Y_COORD_19_112_2: value  <=  8;
            Y_COORD_19_113_0: value  <=  9;
            Y_COORD_19_113_1: value  <=  10;
            Y_COORD_19_114_0: value  <=  7;
            Y_COORD_19_114_1: value  <=  8;
            Y_COORD_19_115_0: value  <=  2;
            Y_COORD_19_115_1: value  <=  5;
            Y_COORD_19_116_0: value  <=  9;
            Y_COORD_19_116_1: value  <=  9;
            Y_COORD_19_117_0: value  <=  9;
            Y_COORD_19_117_1: value  <=  10;
            Y_COORD_19_118_0: value  <=  2;
            Y_COORD_19_118_1: value  <=  5;
            Y_COORD_19_119_0: value  <=  3;
            Y_COORD_19_119_1: value  <=  3;
            Y_COORD_19_120_0: value  <=  3;
            Y_COORD_19_120_1: value  <=  3;
            Y_COORD_19_121_0: value  <=  14;
            Y_COORD_19_121_1: value  <=  15;
            Y_COORD_19_122_0: value  <=  9;
            Y_COORD_19_122_1: value  <=  9;
            Y_COORD_19_123_0: value  <=  9;
            Y_COORD_19_123_1: value  <=  10;
            Y_COORD_19_124_0: value  <=  9;
            Y_COORD_19_124_1: value  <=  10;
            Y_COORD_19_125_0: value  <=  5;
            Y_COORD_19_125_1: value  <=  5;
            Y_COORD_19_125_2: value  <=  9;
            Y_COORD_19_126_0: value  <=  5;
            Y_COORD_19_126_1: value  <=  5;
            Y_COORD_19_126_2: value  <=  9;
            Y_COORD_19_127_0: value  <=  1;
            Y_COORD_19_127_1: value  <=  4;
            Y_COORD_19_128_0: value  <=  0;
            Y_COORD_19_128_1: value  <=  0;
            Y_COORD_19_129_0: value  <=  11;
            Y_COORD_19_129_1: value  <=  11;
            Y_COORD_19_130_0: value  <=  11;
            Y_COORD_19_130_1: value  <=  11;
            Y_COORD_19_131_0: value  <=  4;
            Y_COORD_19_131_1: value  <=  4;
            Y_COORD_19_132_0: value  <=  0;
            Y_COORD_19_132_1: value  <=  0;
            Y_COORD_19_133_0: value  <=  0;
            Y_COORD_19_133_1: value  <=  0;
            Y_COORD_19_134_0: value  <=  1;
            Y_COORD_19_134_1: value  <=  1;
            Y_COORD_19_135_0: value  <=  0;
            Y_COORD_19_135_1: value  <=  0;
            Y_COORD_19_136_0: value  <=  11;
            Y_COORD_19_136_1: value  <=  11;
            Y_COORD_19_137_0: value  <=  0;
            Y_COORD_19_137_1: value  <=  0;
            Y_COORD_19_138_0: value  <=  4;
            Y_COORD_19_138_1: value  <=  4;
            Y_COORD_19_139_0: value  <=  7;
            Y_COORD_19_139_1: value  <=  8;
            Y_COORD_19_140_0: value  <=  1;
            Y_COORD_19_140_1: value  <=  4;
            Y_COORD_19_141_0: value  <=  7;
            Y_COORD_19_141_1: value  <=  8;
            Y_COORD_19_142_0: value  <=  16;
            Y_COORD_19_142_1: value  <=  17;
            Y_COORD_19_143_0: value  <=  8;
            Y_COORD_19_143_1: value  <=  8;
            Y_COORD_19_143_2: value  <=  13;
            Y_COORD_19_144_0: value  <=  9;
            Y_COORD_19_144_1: value  <=  10;
            Y_COORD_19_145_0: value  <=  11;
            Y_COORD_19_145_1: value  <=  11;
            Y_COORD_19_145_2: value  <=  12;
            Y_COORD_19_146_0: value  <=  15;
            Y_COORD_19_146_1: value  <=  16;
            Y_COORD_19_147_0: value  <=  7;
            Y_COORD_19_147_1: value  <=  8;
            Y_COORD_19_148_0: value  <=  7;
            Y_COORD_19_148_1: value  <=  8;
            Y_COORD_19_149_0: value  <=  5;
            Y_COORD_19_149_1: value  <=  8;
            Y_COORD_19_150_0: value  <=  0;
            Y_COORD_19_150_1: value  <=  0;
            Y_COORD_19_151_0: value  <=  2;
            Y_COORD_19_151_1: value  <=  2;
            Y_COORD_19_152_0: value  <=  11;
            Y_COORD_19_152_1: value  <=  11;
            Y_COORD_19_152_2: value  <=  12;
            Y_COORD_19_153_0: value  <=  15;
            Y_COORD_19_153_1: value  <=  16;
            Y_COORD_19_154_0: value  <=  15;
            Y_COORD_19_154_1: value  <=  16;
            Y_COORD_19_155_0: value  <=  12;
            Y_COORD_19_155_1: value  <=  12;
            Y_COORD_19_155_2: value  <=  16;
            Y_COORD_19_156_0: value  <=  8;
            Y_COORD_19_156_1: value  <=  8;
            Y_COORD_19_157_0: value  <=  2;
            Y_COORD_19_157_1: value  <=  2;
            Y_COORD_19_158_0: value  <=  1;
            Y_COORD_19_158_1: value  <=  1;
            Y_COORD_19_159_0: value  <=  2;
            Y_COORD_19_159_1: value  <=  2;
            Y_COORD_19_160_0: value  <=  2;
            Y_COORD_19_160_1: value  <=  2;
            Y_COORD_19_161_0: value  <=  9;
            Y_COORD_19_161_1: value  <=  9;
            Y_COORD_19_161_2: value  <=  11;
            Y_COORD_19_162_0: value  <=  15;
            Y_COORD_19_162_1: value  <=  15;
            Y_COORD_19_162_2: value  <=  16;
            Y_COORD_19_163_0: value  <=  14;
            Y_COORD_19_163_1: value  <=  15;
            Y_COORD_19_164_0: value  <=  13;
            Y_COORD_19_164_1: value  <=  13;
            Y_COORD_19_164_2: value  <=  14;
            Y_COORD_19_165_0: value  <=  9;
            Y_COORD_19_165_1: value  <=  9;
            Y_COORD_19_165_2: value  <=  13;
            Y_COORD_19_166_0: value  <=  13;
            Y_COORD_19_166_1: value  <=  16;
            Y_COORD_19_167_0: value  <=  12;
            Y_COORD_19_167_1: value  <=  13;
            Y_COORD_19_168_0: value  <=  12;
            Y_COORD_19_168_1: value  <=  12;
            Y_COORD_19_168_2: value  <=  13;
            Y_COORD_19_169_0: value  <=  11;
            Y_COORD_19_169_1: value  <=  11;
            Y_COORD_19_169_2: value  <=  13;
            Y_COORD_19_170_0: value  <=  5;
            Y_COORD_19_170_1: value  <=  6;
            Y_COORD_19_171_0: value  <=  10;
            Y_COORD_19_171_1: value  <=  10;
            Y_COORD_19_172_0: value  <=  14;
            Y_COORD_19_172_1: value  <=  15;
            Y_COORD_19_173_0: value  <=  8;
            Y_COORD_19_173_1: value  <=  8;
            Y_COORD_19_173_2: value  <=  14;
            Y_COORD_19_174_0: value  <=  8;
            Y_COORD_19_174_1: value  <=  8;
            Y_COORD_19_174_2: value  <=  14;
            Y_COORD_19_175_0: value  <=  0;
            Y_COORD_19_175_1: value  <=  0;
            Y_COORD_19_176_0: value  <=  11;
            Y_COORD_19_176_1: value  <=  11;
            Y_COORD_19_176_2: value  <=  13;
            Y_COORD_19_177_0: value  <=  16;
            Y_COORD_19_177_1: value  <=  16;
            Y_COORD_19_177_2: value  <=  18;
            Y_COORD_19_178_0: value  <=  7;
            Y_COORD_19_178_1: value  <=  7;
            Y_COORD_19_179_0: value  <=  2;
            Y_COORD_19_179_1: value  <=  2;
            Y_COORD_19_180_0: value  <=  1;
            Y_COORD_19_180_1: value  <=  1;
            Y_COORD_19_181_0: value  <=  19;
            Y_COORD_19_181_1: value  <=  19;
            Y_COORD_20_0_0: value  <=  2;
            Y_COORD_20_0_1: value  <=  2;
            Y_COORD_20_1_0: value  <=  5;
            Y_COORD_20_1_1: value  <=  5;
            Y_COORD_20_2_0: value  <=  4;
            Y_COORD_20_2_1: value  <=  6;
            Y_COORD_20_3_0: value  <=  5;
            Y_COORD_20_3_1: value  <=  9;
            Y_COORD_20_4_0: value  <=  6;
            Y_COORD_20_4_1: value  <=  12;
            Y_COORD_20_5_0: value  <=  6;
            Y_COORD_20_5_1: value  <=  9;
            Y_COORD_20_6_0: value  <=  6;
            Y_COORD_20_6_1: value  <=  9;
            Y_COORD_20_7_0: value  <=  15;
            Y_COORD_20_7_1: value  <=  15;
            Y_COORD_20_7_2: value  <=  17;
            Y_COORD_20_8_0: value  <=  18;
            Y_COORD_20_8_1: value  <=  18;
            Y_COORD_20_9_0: value  <=  3;
            Y_COORD_20_9_1: value  <=  4;
            Y_COORD_20_10_0: value  <=  0;
            Y_COORD_20_10_1: value  <=  2;
            Y_COORD_20_11_0: value  <=  3;
            Y_COORD_20_11_1: value  <=  4;
            Y_COORD_20_12_0: value  <=  11;
            Y_COORD_20_12_1: value  <=  12;
            Y_COORD_20_13_0: value  <=  3;
            Y_COORD_20_13_1: value  <=  4;
            Y_COORD_20_14_0: value  <=  3;
            Y_COORD_20_14_1: value  <=  4;
            Y_COORD_20_15_0: value  <=  0;
            Y_COORD_20_15_1: value  <=  0;
            Y_COORD_20_16_0: value  <=  14;
            Y_COORD_20_16_1: value  <=  16;
            Y_COORD_20_17_0: value  <=  16;
            Y_COORD_20_17_1: value  <=  17;
            Y_COORD_20_18_0: value  <=  6;
            Y_COORD_20_18_1: value  <=  6;
            Y_COORD_20_19_0: value  <=  11;
            Y_COORD_20_19_1: value  <=  12;
            Y_COORD_20_20_0: value  <=  5;
            Y_COORD_20_20_1: value  <=  6;
            Y_COORD_20_21_0: value  <=  9;
            Y_COORD_20_21_1: value  <=  10;
            Y_COORD_20_22_0: value  <=  1;
            Y_COORD_20_22_1: value  <=  1;
            Y_COORD_20_23_0: value  <=  0;
            Y_COORD_20_23_1: value  <=  0;
            Y_COORD_20_24_0: value  <=  0;
            Y_COORD_20_24_1: value  <=  0;
            Y_COORD_20_25_0: value  <=  11;
            Y_COORD_20_25_1: value  <=  12;
            Y_COORD_20_26_0: value  <=  4;
            Y_COORD_20_26_1: value  <=  4;
            Y_COORD_20_27_0: value  <=  3;
            Y_COORD_20_27_1: value  <=  5;
            Y_COORD_20_28_0: value  <=  3;
            Y_COORD_20_28_1: value  <=  5;
            Y_COORD_20_29_0: value  <=  2;
            Y_COORD_20_29_1: value  <=  2;
            Y_COORD_20_29_2: value  <=  5;
            Y_COORD_20_30_0: value  <=  10;
            Y_COORD_20_30_1: value  <=  11;
            Y_COORD_20_31_0: value  <=  2;
            Y_COORD_20_31_1: value  <=  2;
            Y_COORD_20_31_2: value  <=  5;
            Y_COORD_20_32_0: value  <=  11;
            Y_COORD_20_32_1: value  <=  12;
            Y_COORD_20_33_0: value  <=  13;
            Y_COORD_20_33_1: value  <=  14;
            Y_COORD_20_34_0: value  <=  12;
            Y_COORD_20_34_1: value  <=  13;
            Y_COORD_20_35_0: value  <=  11;
            Y_COORD_20_35_1: value  <=  12;
            Y_COORD_20_36_0: value  <=  13;
            Y_COORD_20_36_1: value  <=  14;
            Y_COORD_20_37_0: value  <=  12;
            Y_COORD_20_37_1: value  <=  13;
            Y_COORD_20_38_0: value  <=  11;
            Y_COORD_20_38_1: value  <=  13;
            Y_COORD_20_39_0: value  <=  4;
            Y_COORD_20_39_1: value  <=  4;
            Y_COORD_20_40_0: value  <=  4;
            Y_COORD_20_40_1: value  <=  4;
            Y_COORD_20_41_0: value  <=  5;
            Y_COORD_20_41_1: value  <=  5;
            Y_COORD_20_42_0: value  <=  6;
            Y_COORD_20_42_1: value  <=  6;
            Y_COORD_20_43_0: value  <=  5;
            Y_COORD_20_43_1: value  <=  5;
            Y_COORD_20_44_0: value  <=  13;
            Y_COORD_20_44_1: value  <=  14;
            Y_COORD_20_45_0: value  <=  5;
            Y_COORD_20_45_1: value  <=  5;
            Y_COORD_20_46_0: value  <=  5;
            Y_COORD_20_46_1: value  <=  5;
            Y_COORD_20_47_0: value  <=  9;
            Y_COORD_20_47_1: value  <=  9;
            Y_COORD_20_48_0: value  <=  9;
            Y_COORD_20_48_1: value  <=  9;
            Y_COORD_20_49_0: value  <=  11;
            Y_COORD_20_49_1: value  <=  12;
            Y_COORD_20_50_0: value  <=  11;
            Y_COORD_20_50_1: value  <=  12;
            Y_COORD_20_51_0: value  <=  13;
            Y_COORD_20_51_1: value  <=  14;
            Y_COORD_20_52_0: value  <=  10;
            Y_COORD_20_52_1: value  <=  10;
            Y_COORD_20_52_2: value  <=  12;
            Y_COORD_20_53_0: value  <=  3;
            Y_COORD_20_53_1: value  <=  3;
            Y_COORD_20_54_0: value  <=  2;
            Y_COORD_20_54_1: value  <=  2;
            Y_COORD_20_55_0: value  <=  12;
            Y_COORD_20_55_1: value  <=  12;
            Y_COORD_20_55_2: value  <=  15;
            Y_COORD_20_56_0: value  <=  7;
            Y_COORD_20_56_1: value  <=  7;
            Y_COORD_20_57_0: value  <=  4;
            Y_COORD_20_57_1: value  <=  5;
            Y_COORD_20_58_0: value  <=  7;
            Y_COORD_20_58_1: value  <=  7;
            Y_COORD_20_59_0: value  <=  2;
            Y_COORD_20_59_1: value  <=  4;
            Y_COORD_20_60_0: value  <=  16;
            Y_COORD_20_60_1: value  <=  16;
            Y_COORD_20_61_0: value  <=  13;
            Y_COORD_20_61_1: value  <=  14;
            Y_COORD_20_62_0: value  <=  7;
            Y_COORD_20_62_1: value  <=  7;
            Y_COORD_20_63_0: value  <=  10;
            Y_COORD_20_63_1: value  <=  12;
            Y_COORD_20_64_0: value  <=  10;
            Y_COORD_20_64_1: value  <=  10;
            Y_COORD_20_65_0: value  <=  9;
            Y_COORD_20_65_1: value  <=  10;
            Y_COORD_20_66_0: value  <=  9;
            Y_COORD_20_66_1: value  <=  10;
            Y_COORD_20_67_0: value  <=  7;
            Y_COORD_20_67_1: value  <=  7;
            Y_COORD_20_67_2: value  <=  8;
            Y_COORD_20_68_0: value  <=  7;
            Y_COORD_20_68_1: value  <=  7;
            Y_COORD_20_68_2: value  <=  8;
            Y_COORD_20_69_0: value  <=  0;
            Y_COORD_20_69_1: value  <=  0;
            Y_COORD_20_70_0: value  <=  0;
            Y_COORD_20_70_1: value  <=  0;
            Y_COORD_20_71_0: value  <=  4;
            Y_COORD_20_71_1: value  <=  4;
            Y_COORD_20_72_0: value  <=  14;
            Y_COORD_20_72_1: value  <=  15;
            Y_COORD_20_73_0: value  <=  14;
            Y_COORD_20_73_1: value  <=  15;
            Y_COORD_20_74_0: value  <=  2;
            Y_COORD_20_74_1: value  <=  2;
            Y_COORD_20_75_0: value  <=  2;
            Y_COORD_20_75_1: value  <=  7;
            Y_COORD_20_76_0: value  <=  14;
            Y_COORD_20_76_1: value  <=  15;
            Y_COORD_20_77_0: value  <=  2;
            Y_COORD_20_77_1: value  <=  2;
            Y_COORD_20_77_2: value  <=  8;
            Y_COORD_20_78_0: value  <=  7;
            Y_COORD_20_78_1: value  <=  8;
            Y_COORD_20_79_0: value  <=  13;
            Y_COORD_20_79_1: value  <=  16;
            Y_COORD_20_80_0: value  <=  6;
            Y_COORD_20_80_1: value  <=  7;
            Y_COORD_20_81_0: value  <=  2;
            Y_COORD_20_81_1: value  <=  4;
            Y_COORD_20_82_0: value  <=  6;
            Y_COORD_20_82_1: value  <=  6;
            Y_COORD_20_82_2: value  <=  7;
            Y_COORD_20_83_0: value  <=  2;
            Y_COORD_20_83_1: value  <=  4;
            Y_COORD_20_84_0: value  <=  2;
            Y_COORD_20_84_1: value  <=  4;
            Y_COORD_20_85_0: value  <=  6;
            Y_COORD_20_85_1: value  <=  6;
            Y_COORD_20_86_0: value  <=  4;
            Y_COORD_20_86_1: value  <=  9;
            Y_COORD_20_87_0: value  <=  5;
            Y_COORD_20_87_1: value  <=  5;
            Y_COORD_20_88_0: value  <=  13;
            Y_COORD_20_88_1: value  <=  14;
            Y_COORD_20_89_0: value  <=  13;
            Y_COORD_20_89_1: value  <=  14;
            Y_COORD_20_90_0: value  <=  16;
            Y_COORD_20_90_1: value  <=  16;
            Y_COORD_20_90_2: value  <=  18;
            Y_COORD_20_91_0: value  <=  6;
            Y_COORD_20_91_1: value  <=  6;
            Y_COORD_20_91_2: value  <=  9;
            Y_COORD_20_92_0: value  <=  14;
            Y_COORD_20_92_1: value  <=  15;
            Y_COORD_20_93_0: value  <=  16;
            Y_COORD_20_93_1: value  <=  17;
            Y_COORD_20_94_0: value  <=  4;
            Y_COORD_20_94_1: value  <=  5;
            Y_COORD_20_95_0: value  <=  4;
            Y_COORD_20_95_1: value  <=  5;
            Y_COORD_20_96_0: value  <=  4;
            Y_COORD_20_96_1: value  <=  6;
            Y_COORD_20_97_0: value  <=  11;
            Y_COORD_20_97_1: value  <=  14;
            Y_COORD_20_98_0: value  <=  11;
            Y_COORD_20_98_1: value  <=  14;
            Y_COORD_20_99_0: value  <=  7;
            Y_COORD_20_99_1: value  <=  7;
            Y_COORD_20_100_0: value  <=  0;
            Y_COORD_20_100_1: value  <=  0;
            Y_COORD_20_101_0: value  <=  3;
            Y_COORD_20_101_1: value  <=  3;
            Y_COORD_20_102_0: value  <=  2;
            Y_COORD_20_102_1: value  <=  2;
            Y_COORD_20_103_0: value  <=  2;
            Y_COORD_20_103_1: value  <=  2;
            Y_COORD_20_103_2: value  <=  3;
            Y_COORD_20_104_0: value  <=  1;
            Y_COORD_20_104_1: value  <=  3;
            Y_COORD_20_105_0: value  <=  17;
            Y_COORD_20_105_1: value  <=  18;
            Y_COORD_20_106_0: value  <=  0;
            Y_COORD_20_106_1: value  <=  0;
            Y_COORD_20_107_0: value  <=  0;
            Y_COORD_20_107_1: value  <=  1;
            Y_COORD_20_108_0: value  <=  14;
            Y_COORD_20_108_1: value  <=  15;
            Y_COORD_20_109_0: value  <=  12;
            Y_COORD_20_109_1: value  <=  12;
            Y_COORD_20_109_2: value  <=  16;
            Y_COORD_20_110_0: value  <=  0;
            Y_COORD_20_110_1: value  <=  1;
            Y_COORD_20_111_0: value  <=  12;
            Y_COORD_20_111_1: value  <=  12;
            Y_COORD_20_111_2: value  <=  16;
            Y_COORD_20_112_0: value  <=  0;
            Y_COORD_20_112_1: value  <=  0;
            Y_COORD_20_112_2: value  <=  6;
            Y_COORD_20_113_0: value  <=  1;
            Y_COORD_20_113_1: value  <=  4;
            Y_COORD_20_114_0: value  <=  2;
            Y_COORD_20_114_1: value  <=  3;
            Y_COORD_20_115_0: value  <=  14;
            Y_COORD_20_115_1: value  <=  14;
            Y_COORD_20_115_2: value  <=  17;
            Y_COORD_20_116_0: value  <=  17;
            Y_COORD_20_116_1: value  <=  17;
            Y_COORD_20_116_2: value  <=  18;
            Y_COORD_20_117_0: value  <=  3;
            Y_COORD_20_117_1: value  <=  3;
            Y_COORD_20_117_2: value  <=  6;
            Y_COORD_20_118_0: value  <=  12;
            Y_COORD_20_118_1: value  <=  12;
            Y_COORD_20_119_0: value  <=  7;
            Y_COORD_20_119_1: value  <=  7;
            Y_COORD_20_120_0: value  <=  15;
            Y_COORD_20_120_1: value  <=  15;
            Y_COORD_20_121_0: value  <=  4;
            Y_COORD_20_121_1: value  <=  4;
            Y_COORD_20_122_0: value  <=  7;
            Y_COORD_20_122_1: value  <=  7;
            Y_COORD_20_123_0: value  <=  3;
            Y_COORD_20_123_1: value  <=  3;
            Y_COORD_20_124_0: value  <=  3;
            Y_COORD_20_124_1: value  <=  3;
            Y_COORD_20_125_0: value  <=  7;
            Y_COORD_20_125_1: value  <=  7;
            Y_COORD_20_126_0: value  <=  17;
            Y_COORD_20_126_1: value  <=  17;
            Y_COORD_20_127_0: value  <=  14;
            Y_COORD_20_127_1: value  <=  14;
            Y_COORD_20_127_2: value  <=  17;
            Y_COORD_20_128_0: value  <=  13;
            Y_COORD_20_128_1: value  <=  13;
            Y_COORD_20_128_2: value  <=  15;
            Y_COORD_20_129_0: value  <=  5;
            Y_COORD_20_129_1: value  <=  5;
            Y_COORD_20_129_2: value  <=  6;
            Y_COORD_20_130_0: value  <=  2;
            Y_COORD_20_130_1: value  <=  2;
            Y_COORD_20_130_2: value  <=  8;
            Y_COORD_20_131_0: value  <=  1;
            Y_COORD_20_131_1: value  <=  2;
            Y_COORD_20_132_0: value  <=  16;
            Y_COORD_20_132_1: value  <=  17;
            Y_COORD_20_133_0: value  <=  17;
            Y_COORD_20_133_1: value  <=  17;
            Y_COORD_20_134_0: value  <=  15;
            Y_COORD_20_134_1: value  <=  15;
            Y_COORD_20_134_2: value  <=  16;
            Y_COORD_20_135_0: value  <=  15;
            Y_COORD_20_135_1: value  <=  16;
            Y_COORD_20_136_0: value  <=  16;
            Y_COORD_20_136_1: value  <=  16;
            Y_COORD_20_136_2: value  <=  18;
            Y_COORD_20_137_0: value  <=  11;
            Y_COORD_20_137_1: value  <=  14;
            Y_COORD_20_138_0: value  <=  13;
            Y_COORD_20_138_1: value  <=  14;
            Y_COORD_20_139_0: value  <=  14;
            Y_COORD_20_139_1: value  <=  14;
            Y_COORD_20_139_2: value  <=  17;
            Y_COORD_20_140_0: value  <=  9;
            Y_COORD_20_140_1: value  <=  9;
            Y_COORD_20_141_0: value  <=  14;
            Y_COORD_20_141_1: value  <=  14;
            Y_COORD_20_141_2: value  <=  17;
            Y_COORD_20_142_0: value  <=  2;
            Y_COORD_20_142_1: value  <=  4;
            Y_COORD_20_143_0: value  <=  0;
            Y_COORD_20_143_1: value  <=  10;
            Y_COORD_20_144_0: value  <=  14;
            Y_COORD_20_144_1: value  <=  14;
            Y_COORD_20_144_2: value  <=  17;
            Y_COORD_20_145_0: value  <=  14;
            Y_COORD_20_145_1: value  <=  14;
            Y_COORD_20_145_2: value  <=  17;
            Y_COORD_20_146_0: value  <=  11;
            Y_COORD_20_146_1: value  <=  11;
            Y_COORD_20_147_0: value  <=  17;
            Y_COORD_20_147_1: value  <=  17;
            Y_COORD_20_148_0: value  <=  17;
            Y_COORD_20_148_1: value  <=  17;
            Y_COORD_20_149_0: value  <=  14;
            Y_COORD_20_149_1: value  <=  14;
            Y_COORD_20_149_2: value  <=  17;
            Y_COORD_20_150_0: value  <=  14;
            Y_COORD_20_150_1: value  <=  14;
            Y_COORD_20_150_2: value  <=  17;
            Y_COORD_20_151_0: value  <=  14;
            Y_COORD_20_151_1: value  <=  14;
            Y_COORD_20_151_2: value  <=  17;
            Y_COORD_20_152_0: value  <=  14;
            Y_COORD_20_152_1: value  <=  14;
            Y_COORD_20_152_2: value  <=  17;
            Y_COORD_20_153_0: value  <=  0;
            Y_COORD_20_153_1: value  <=  4;
            Y_COORD_20_154_0: value  <=  7;
            Y_COORD_20_154_1: value  <=  7;
            Y_COORD_20_155_0: value  <=  3;
            Y_COORD_20_155_1: value  <=  3;
            Y_COORD_20_156_0: value  <=  3;
            Y_COORD_20_156_1: value  <=  3;
            Y_COORD_20_157_0: value  <=  8;
            Y_COORD_20_157_1: value  <=  9;
            Y_COORD_20_158_0: value  <=  11;
            Y_COORD_20_158_1: value  <=  11;
            Y_COORD_20_159_0: value  <=  12;
            Y_COORD_20_159_1: value  <=  12;
            Y_COORD_20_159_2: value  <=  16;
            Y_COORD_20_160_0: value  <=  6;
            Y_COORD_20_160_1: value  <=  6;
            Y_COORD_20_161_0: value  <=  11;
            Y_COORD_20_161_1: value  <=  11;
            Y_COORD_20_162_0: value  <=  13;
            Y_COORD_20_162_1: value  <=  13;
            Y_COORD_20_163_0: value  <=  9;
            Y_COORD_20_163_1: value  <=  10;
            Y_COORD_20_164_0: value  <=  3;
            Y_COORD_20_164_1: value  <=  4;
            Y_COORD_20_165_0: value  <=  3;
            Y_COORD_20_165_1: value  <=  4;
            Y_COORD_20_166_0: value  <=  4;
            Y_COORD_20_166_1: value  <=  8;
            Y_COORD_20_167_0: value  <=  3;
            Y_COORD_20_167_1: value  <=  4;
            Y_COORD_20_168_0: value  <=  8;
            Y_COORD_20_168_1: value  <=  9;
            Y_COORD_20_169_0: value  <=  3;
            Y_COORD_20_169_1: value  <=  4;
            Y_COORD_20_170_0: value  <=  11;
            Y_COORD_20_170_1: value  <=  11;
            Y_COORD_20_171_0: value  <=  12;
            Y_COORD_20_171_1: value  <=  12;
            Y_COORD_20_171_2: value  <=  16;
            Y_COORD_20_172_0: value  <=  8;
            Y_COORD_20_172_1: value  <=  9;
            Y_COORD_20_173_0: value  <=  13;
            Y_COORD_20_173_1: value  <=  13;
            Y_COORD_20_173_2: value  <=  14;
            Y_COORD_20_174_0: value  <=  13;
            Y_COORD_20_174_1: value  <=  14;
            Y_COORD_20_175_0: value  <=  12;
            Y_COORD_20_175_1: value  <=  12;
            Y_COORD_20_176_0: value  <=  3;
            Y_COORD_20_176_1: value  <=  4;
            Y_COORD_20_177_0: value  <=  4;
            Y_COORD_20_177_1: value  <=  5;
            Y_COORD_20_178_0: value  <=  2;
            Y_COORD_20_178_1: value  <=  3;
            Y_COORD_20_179_0: value  <=  12;
            Y_COORD_20_179_1: value  <=  12;
            Y_COORD_20_179_2: value  <=  16;
            Y_COORD_20_180_0: value  <=  12;
            Y_COORD_20_180_1: value  <=  12;
            Y_COORD_20_180_2: value  <=  16;
            Y_COORD_20_181_0: value  <=  13;
            Y_COORD_20_181_1: value  <=  15;
            Y_COORD_20_182_0: value  <=  13;
            Y_COORD_20_182_1: value  <=  15;
            Y_COORD_20_183_0: value  <=  5;
            Y_COORD_20_183_1: value  <=  5;
            Y_COORD_20_183_2: value  <=  6;
            Y_COORD_20_184_0: value  <=  14;
            Y_COORD_20_184_1: value  <=  17;
            Y_COORD_20_185_0: value  <=  14;
            Y_COORD_20_185_1: value  <=  15;
            Y_COORD_20_186_0: value  <=  16;
            Y_COORD_20_186_1: value  <=  16;
            Y_COORD_20_186_2: value  <=  17;
            Y_COORD_20_187_0: value  <=  6;
            Y_COORD_20_187_1: value  <=  7;
            Y_COORD_20_188_0: value  <=  17;
            Y_COORD_20_188_1: value  <=  17;
            Y_COORD_20_188_2: value  <=  18;
            Y_COORD_20_189_0: value  <=  6;
            Y_COORD_20_189_1: value  <=  7;
            Y_COORD_20_190_0: value  <=  13;
            Y_COORD_20_190_1: value  <=  13;
            Y_COORD_20_191_0: value  <=  2;
            Y_COORD_20_191_1: value  <=  2;
            Y_COORD_20_192_0: value  <=  18;
            Y_COORD_20_192_1: value  <=  18;
            Y_COORD_20_192_2: value  <=  19;
            Y_COORD_20_193_0: value  <=  16;
            Y_COORD_20_193_1: value  <=  16;
            Y_COORD_20_194_0: value  <=  6;
            Y_COORD_20_194_1: value  <=  7;
            Y_COORD_20_195_0: value  <=  1;
            Y_COORD_20_195_1: value  <=  2;
            Y_COORD_20_196_0: value  <=  14;
            Y_COORD_20_196_1: value  <=  14;
            Y_COORD_20_196_2: value  <=  15;
            Y_COORD_20_197_0: value  <=  3;
            Y_COORD_20_197_1: value  <=  3;
            Y_COORD_20_198_0: value  <=  13;
            Y_COORD_20_198_1: value  <=  13;
            Y_COORD_20_199_0: value  <=  11;
            Y_COORD_20_199_1: value  <=  12;
            Y_COORD_20_200_0: value  <=  15;
            Y_COORD_20_200_1: value  <=  15;
            Y_COORD_20_200_2: value  <=  17;
            Y_COORD_20_201_0: value  <=  7;
            Y_COORD_20_201_1: value  <=  7;
            Y_COORD_20_201_2: value  <=  8;
            Y_COORD_20_202_0: value  <=  11;
            Y_COORD_20_202_1: value  <=  12;
            Y_COORD_20_203_0: value  <=  0;
            Y_COORD_20_203_1: value  <=  0;
            Y_COORD_20_204_0: value  <=  11;
            Y_COORD_20_204_1: value  <=  12;
            Y_COORD_20_205_0: value  <=  0;
            Y_COORD_20_205_1: value  <=  0;
            Y_COORD_20_206_0: value  <=  10;
            Y_COORD_20_206_1: value  <=  10;
            Y_COORD_20_207_0: value  <=  12;
            Y_COORD_20_207_1: value  <=  13;
            Y_COORD_20_208_0: value  <=  6;
            Y_COORD_20_208_1: value  <=  6;
            Y_COORD_20_209_0: value  <=  4;
            Y_COORD_20_209_1: value  <=  4;
            Y_COORD_20_210_0: value  <=  0;
            Y_COORD_20_210_1: value  <=  1;
            Y_COORD_21_0_0: value  <=  3;
            Y_COORD_21_0_1: value  <=  6;
            Y_COORD_21_1_0: value  <=  2;
            Y_COORD_21_1_1: value  <=  2;
            Y_COORD_21_2_0: value  <=  2;
            Y_COORD_21_2_1: value  <=  2;
            Y_COORD_21_3_0: value  <=  4;
            Y_COORD_21_3_1: value  <=  4;
            Y_COORD_21_4_0: value  <=  4;
            Y_COORD_21_4_1: value  <=  4;
            Y_COORD_21_5_0: value  <=  10;
            Y_COORD_21_5_1: value  <=  12;
            Y_COORD_21_6_0: value  <=  10;
            Y_COORD_21_6_1: value  <=  10;
            Y_COORD_21_7_0: value  <=  9;
            Y_COORD_21_7_1: value  <=  12;
            Y_COORD_21_8_0: value  <=  17;
            Y_COORD_21_8_1: value  <=  18;
            Y_COORD_21_9_0: value  <=  3;
            Y_COORD_21_9_1: value  <=  3;
            Y_COORD_21_9_2: value  <=  11;
            Y_COORD_21_10_0: value  <=  9;
            Y_COORD_21_10_1: value  <=  12;
            Y_COORD_21_11_0: value  <=  1;
            Y_COORD_21_11_1: value  <=  2;
            Y_COORD_21_12_0: value  <=  18;
            Y_COORD_21_12_1: value  <=  18;
            Y_COORD_21_12_2: value  <=  19;
            Y_COORD_21_13_0: value  <=  4;
            Y_COORD_21_13_1: value  <=  4;
            Y_COORD_21_13_2: value  <=  9;
            Y_COORD_21_14_0: value  <=  5;
            Y_COORD_21_14_1: value  <=  10;
            Y_COORD_21_15_0: value  <=  8;
            Y_COORD_21_15_1: value  <=  8;
            Y_COORD_21_16_0: value  <=  8;
            Y_COORD_21_16_1: value  <=  8;
            Y_COORD_21_17_0: value  <=  5;
            Y_COORD_21_17_1: value  <=  7;
            Y_COORD_21_18_0: value  <=  7;
            Y_COORD_21_18_1: value  <=  7;
            Y_COORD_21_19_0: value  <=  11;
            Y_COORD_21_19_1: value  <=  12;
            Y_COORD_21_20_0: value  <=  0;
            Y_COORD_21_20_1: value  <=  1;
            Y_COORD_21_21_0: value  <=  2;
            Y_COORD_21_21_1: value  <=  3;
            Y_COORD_21_22_0: value  <=  1;
            Y_COORD_21_22_1: value  <=  7;
            Y_COORD_21_23_0: value  <=  4;
            Y_COORD_21_23_1: value  <=  4;
            Y_COORD_21_24_0: value  <=  13;
            Y_COORD_21_24_1: value  <=  14;
            Y_COORD_21_25_0: value  <=  14;
            Y_COORD_21_25_1: value  <=  16;
            Y_COORD_21_26_0: value  <=  2;
            Y_COORD_21_26_1: value  <=  2;
            Y_COORD_21_27_0: value  <=  1;
            Y_COORD_21_27_1: value  <=  2;
            Y_COORD_21_28_0: value  <=  1;
            Y_COORD_21_28_1: value  <=  2;
            Y_COORD_21_29_0: value  <=  13;
            Y_COORD_21_29_1: value  <=  14;
            Y_COORD_21_30_0: value  <=  13;
            Y_COORD_21_30_1: value  <=  14;
            Y_COORD_21_31_0: value  <=  12;
            Y_COORD_21_31_1: value  <=  13;
            Y_COORD_21_32_0: value  <=  2;
            Y_COORD_21_32_1: value  <=  3;
            Y_COORD_21_33_0: value  <=  6;
            Y_COORD_21_33_1: value  <=  6;
            Y_COORD_21_33_2: value  <=  8;
            Y_COORD_21_34_0: value  <=  13;
            Y_COORD_21_34_1: value  <=  16;
            Y_COORD_21_35_0: value  <=  12;
            Y_COORD_21_35_1: value  <=  12;
            Y_COORD_21_35_2: value  <=  13;
            Y_COORD_21_36_0: value  <=  12;
            Y_COORD_21_36_1: value  <=  13;
            Y_COORD_21_37_0: value  <=  4;
            Y_COORD_21_37_1: value  <=  6;
            Y_COORD_21_38_0: value  <=  17;
            Y_COORD_21_38_1: value  <=  18;
            Y_COORD_21_39_0: value  <=  4;
            Y_COORD_21_39_1: value  <=  6;
            Y_COORD_21_40_0: value  <=  4;
            Y_COORD_21_40_1: value  <=  6;
            Y_COORD_21_41_0: value  <=  6;
            Y_COORD_21_41_1: value  <=  6;
            Y_COORD_21_42_0: value  <=  9;
            Y_COORD_21_42_1: value  <=  9;
            Y_COORD_21_43_0: value  <=  12;
            Y_COORD_21_43_1: value  <=  13;
            Y_COORD_21_44_0: value  <=  12;
            Y_COORD_21_44_1: value  <=  14;
            Y_COORD_21_45_0: value  <=  12;
            Y_COORD_21_45_1: value  <=  13;
            Y_COORD_21_46_0: value  <=  15;
            Y_COORD_21_46_1: value  <=  16;
            Y_COORD_21_47_0: value  <=  9;
            Y_COORD_21_47_1: value  <=  9;
            Y_COORD_21_47_2: value  <=  13;
            Y_COORD_21_48_0: value  <=  12;
            Y_COORD_21_48_1: value  <=  12;
            Y_COORD_21_48_2: value  <=  15;
            Y_COORD_21_49_0: value  <=  11;
            Y_COORD_21_49_1: value  <=  11;
            Y_COORD_21_50_0: value  <=  7;
            Y_COORD_21_50_1: value  <=  7;
            Y_COORD_21_50_2: value  <=  12;
            Y_COORD_21_51_0: value  <=  0;
            Y_COORD_21_51_1: value  <=  0;
            Y_COORD_21_52_0: value  <=  11;
            Y_COORD_21_52_1: value  <=  13;
            Y_COORD_21_53_0: value  <=  12;
            Y_COORD_21_53_1: value  <=  13;
            Y_COORD_21_54_0: value  <=  14;
            Y_COORD_21_54_1: value  <=  14;
            Y_COORD_21_54_2: value  <=  17;
            Y_COORD_21_55_0: value  <=  1;
            Y_COORD_21_55_1: value  <=  1;
            Y_COORD_21_56_0: value  <=  8;
            Y_COORD_21_56_1: value  <=  9;
            Y_COORD_21_57_0: value  <=  9;
            Y_COORD_21_57_1: value  <=  9;
            Y_COORD_21_58_0: value  <=  7;
            Y_COORD_21_58_1: value  <=  8;
            Y_COORD_21_59_0: value  <=  0;
            Y_COORD_21_59_1: value  <=  0;
            Y_COORD_21_60_0: value  <=  0;
            Y_COORD_21_60_1: value  <=  0;
            Y_COORD_21_61_0: value  <=  5;
            Y_COORD_21_61_1: value  <=  5;
            Y_COORD_21_62_0: value  <=  5;
            Y_COORD_21_62_1: value  <=  5;
            Y_COORD_21_63_0: value  <=  0;
            Y_COORD_21_63_1: value  <=  0;
            Y_COORD_21_64_0: value  <=  0;
            Y_COORD_21_64_1: value  <=  0;
            Y_COORD_21_65_0: value  <=  12;
            Y_COORD_21_65_1: value  <=  12;
            Y_COORD_21_65_2: value  <=  13;
            Y_COORD_21_66_0: value  <=  12;
            Y_COORD_21_66_1: value  <=  12;
            Y_COORD_21_66_2: value  <=  13;
            Y_COORD_21_67_0: value  <=  0;
            Y_COORD_21_67_1: value  <=  0;
            Y_COORD_21_68_0: value  <=  11;
            Y_COORD_21_68_1: value  <=  12;
            Y_COORD_21_69_0: value  <=  7;
            Y_COORD_21_69_1: value  <=  8;
            Y_COORD_21_70_0: value  <=  10;
            Y_COORD_21_70_1: value  <=  10;
            Y_COORD_21_71_0: value  <=  9;
            Y_COORD_21_71_1: value  <=  9;
            Y_COORD_21_72_0: value  <=  9;
            Y_COORD_21_72_1: value  <=  9;
            Y_COORD_21_73_0: value  <=  0;
            Y_COORD_21_73_1: value  <=  0;
            Y_COORD_21_74_0: value  <=  0;
            Y_COORD_21_74_1: value  <=  0;
            Y_COORD_21_75_0: value  <=  14;
            Y_COORD_21_75_1: value  <=  14;
            Y_COORD_21_75_2: value  <=  16;
            Y_COORD_21_76_0: value  <=  13;
            Y_COORD_21_76_1: value  <=  14;
            Y_COORD_21_77_0: value  <=  10;
            Y_COORD_21_77_1: value  <=  14;
            Y_COORD_21_78_0: value  <=  10;
            Y_COORD_21_78_1: value  <=  10;
            Y_COORD_21_78_2: value  <=  14;
            Y_COORD_21_79_0: value  <=  8;
            Y_COORD_21_79_1: value  <=  8;
            Y_COORD_21_80_0: value  <=  12;
            Y_COORD_21_80_1: value  <=  15;
            Y_COORD_21_81_0: value  <=  8;
            Y_COORD_21_81_1: value  <=  8;
            Y_COORD_21_82_0: value  <=  8;
            Y_COORD_21_82_1: value  <=  8;
            Y_COORD_21_83_0: value  <=  2;
            Y_COORD_21_83_1: value  <=  9;
            Y_COORD_21_84_0: value  <=  1;
            Y_COORD_21_84_1: value  <=  1;
            Y_COORD_21_84_2: value  <=  6;
            Y_COORD_21_85_0: value  <=  14;
            Y_COORD_21_85_1: value  <=  15;
            Y_COORD_21_86_0: value  <=  7;
            Y_COORD_21_86_1: value  <=  7;
            Y_COORD_21_87_0: value  <=  4;
            Y_COORD_21_87_1: value  <=  5;
            Y_COORD_21_88_0: value  <=  4;
            Y_COORD_21_88_1: value  <=  5;
            Y_COORD_21_89_0: value  <=  5;
            Y_COORD_21_89_1: value  <=  5;
            Y_COORD_21_89_2: value  <=  6;
            Y_COORD_21_90_0: value  <=  19;
            Y_COORD_21_90_1: value  <=  19;
            Y_COORD_21_91_0: value  <=  12;
            Y_COORD_21_91_1: value  <=  14;
            Y_COORD_21_92_0: value  <=  15;
            Y_COORD_21_92_1: value  <=  16;
            Y_COORD_21_93_0: value  <=  16;
            Y_COORD_21_93_1: value  <=  16;
            Y_COORD_21_94_0: value  <=  10;
            Y_COORD_21_94_1: value  <=  10;
            Y_COORD_21_95_0: value  <=  8;
            Y_COORD_21_95_1: value  <=  8;
            Y_COORD_21_96_0: value  <=  8;
            Y_COORD_21_96_1: value  <=  8;
            Y_COORD_21_97_0: value  <=  14;
            Y_COORD_21_97_1: value  <=  14;
            Y_COORD_21_98_0: value  <=  1;
            Y_COORD_21_98_1: value  <=  1;
            Y_COORD_21_99_0: value  <=  7;
            Y_COORD_21_99_1: value  <=  7;
            Y_COORD_21_100_0: value  <=  6;
            Y_COORD_21_100_1: value  <=  6;
            Y_COORD_21_101_0: value  <=  8;
            Y_COORD_21_101_1: value  <=  9;
            Y_COORD_21_102_0: value  <=  11;
            Y_COORD_21_102_1: value  <=  11;
            Y_COORD_21_102_2: value  <=  14;
            Y_COORD_21_103_0: value  <=  7;
            Y_COORD_21_103_1: value  <=  7;
            Y_COORD_21_103_2: value  <=  8;
            Y_COORD_21_104_0: value  <=  5;
            Y_COORD_21_104_1: value  <=  6;
            Y_COORD_21_105_0: value  <=  7;
            Y_COORD_21_105_1: value  <=  7;
            Y_COORD_21_106_0: value  <=  1;
            Y_COORD_21_106_1: value  <=  7;
            Y_COORD_21_107_0: value  <=  5;
            Y_COORD_21_107_1: value  <=  6;
            Y_COORD_21_108_0: value  <=  5;
            Y_COORD_21_108_1: value  <=  6;
            Y_COORD_21_109_0: value  <=  4;
            Y_COORD_21_109_1: value  <=  5;
            Y_COORD_21_110_0: value  <=  14;
            Y_COORD_21_110_1: value  <=  15;
            Y_COORD_21_111_0: value  <=  4;
            Y_COORD_21_111_1: value  <=  5;
            Y_COORD_21_112_0: value  <=  4;
            Y_COORD_21_112_1: value  <=  5;
            Y_COORD_21_113_0: value  <=  14;
            Y_COORD_21_113_1: value  <=  14;
            Y_COORD_21_113_2: value  <=  17;
            Y_COORD_21_114_0: value  <=  14;
            Y_COORD_21_114_1: value  <=  14;
            Y_COORD_21_115_0: value  <=  5;
            Y_COORD_21_115_1: value  <=  5;
            Y_COORD_21_116_0: value  <=  5;
            Y_COORD_21_116_1: value  <=  5;
            Y_COORD_21_117_0: value  <=  13;
            Y_COORD_21_117_1: value  <=  14;
            Y_COORD_21_118_0: value  <=  2;
            Y_COORD_21_118_1: value  <=  3;
            Y_COORD_21_119_0: value  <=  13;
            Y_COORD_21_119_1: value  <=  14;
            Y_COORD_21_120_0: value  <=  7;
            Y_COORD_21_120_1: value  <=  7;
            Y_COORD_21_120_2: value  <=  8;
            Y_COORD_21_121_0: value  <=  5;
            Y_COORD_21_121_1: value  <=  5;
            Y_COORD_21_122_0: value  <=  13;
            Y_COORD_21_122_1: value  <=  14;
            Y_COORD_21_123_0: value  <=  0;
            Y_COORD_21_123_1: value  <=  0;
            Y_COORD_21_124_0: value  <=  3;
            Y_COORD_21_124_1: value  <=  3;
            Y_COORD_21_124_2: value  <=  11;
            Y_COORD_21_125_0: value  <=  0;
            Y_COORD_21_125_1: value  <=  0;
            Y_COORD_21_126_0: value  <=  0;
            Y_COORD_21_126_1: value  <=  0;
            Y_COORD_21_127_0: value  <=  16;
            Y_COORD_21_127_1: value  <=  16;
            Y_COORD_21_128_0: value  <=  16;
            Y_COORD_21_128_1: value  <=  16;
            Y_COORD_21_129_0: value  <=  5;
            Y_COORD_21_129_1: value  <=  5;
            Y_COORD_21_130_0: value  <=  5;
            Y_COORD_21_130_1: value  <=  5;
            Y_COORD_21_131_0: value  <=  6;
            Y_COORD_21_131_1: value  <=  13;
            Y_COORD_21_132_0: value  <=  10;
            Y_COORD_21_132_1: value  <=  12;
            Y_COORD_21_133_0: value  <=  7;
            Y_COORD_21_133_1: value  <=  8;
            Y_COORD_21_134_0: value  <=  1;
            Y_COORD_21_134_1: value  <=  1;
            Y_COORD_21_134_2: value  <=  4;
            Y_COORD_21_135_0: value  <=  7;
            Y_COORD_21_135_1: value  <=  8;
            Y_COORD_21_136_0: value  <=  6;
            Y_COORD_21_136_1: value  <=  13;
            Y_COORD_21_137_0: value  <=  0;
            Y_COORD_21_137_1: value  <=  0;
            Y_COORD_21_138_0: value  <=  6;
            Y_COORD_21_138_1: value  <=  7;
            Y_COORD_21_139_0: value  <=  0;
            Y_COORD_21_139_1: value  <=  8;
            Y_COORD_21_140_0: value  <=  0;
            Y_COORD_21_140_1: value  <=  0;
            Y_COORD_21_141_0: value  <=  0;
            Y_COORD_21_141_1: value  <=  0;
            Y_COORD_21_142_0: value  <=  7;
            Y_COORD_21_142_1: value  <=  8;
            Y_COORD_21_143_0: value  <=  4;
            Y_COORD_21_143_1: value  <=  6;
            Y_COORD_21_144_0: value  <=  7;
            Y_COORD_21_144_1: value  <=  8;
            Y_COORD_21_145_0: value  <=  6;
            Y_COORD_21_145_1: value  <=  9;
            Y_COORD_21_146_0: value  <=  4;
            Y_COORD_21_146_1: value  <=  4;
            Y_COORD_21_147_0: value  <=  0;
            Y_COORD_21_147_1: value  <=  0;
            Y_COORD_21_147_2: value  <=  2;
            Y_COORD_21_148_0: value  <=  2;
            Y_COORD_21_148_1: value  <=  6;
            Y_COORD_21_149_0: value  <=  2;
            Y_COORD_21_149_1: value  <=  6;
            Y_COORD_21_150_0: value  <=  14;
            Y_COORD_21_150_1: value  <=  15;
            Y_COORD_21_151_0: value  <=  14;
            Y_COORD_21_151_1: value  <=  15;
            Y_COORD_21_152_0: value  <=  14;
            Y_COORD_21_152_1: value  <=  15;
            Y_COORD_21_153_0: value  <=  4;
            Y_COORD_21_153_1: value  <=  6;
            Y_COORD_21_154_0: value  <=  4;
            Y_COORD_21_154_1: value  <=  6;
            Y_COORD_21_155_0: value  <=  5;
            Y_COORD_21_155_1: value  <=  6;
            Y_COORD_21_156_0: value  <=  5;
            Y_COORD_21_156_1: value  <=  6;
            Y_COORD_21_157_0: value  <=  0;
            Y_COORD_21_157_1: value  <=  2;
            Y_COORD_21_158_0: value  <=  1;
            Y_COORD_21_158_1: value  <=  1;
            Y_COORD_21_159_0: value  <=  6;
            Y_COORD_21_159_1: value  <=  6;
            Y_COORD_21_160_0: value  <=  5;
            Y_COORD_21_160_1: value  <=  5;
            Y_COORD_21_160_2: value  <=  6;
            Y_COORD_21_161_0: value  <=  5;
            Y_COORD_21_161_1: value  <=  6;
            Y_COORD_21_162_0: value  <=  5;
            Y_COORD_21_162_1: value  <=  6;
            Y_COORD_21_163_0: value  <=  10;
            Y_COORD_21_163_1: value  <=  11;
            Y_COORD_21_164_0: value  <=  8;
            Y_COORD_21_164_1: value  <=  9;
            Y_COORD_21_165_0: value  <=  0;
            Y_COORD_21_165_1: value  <=  3;
            Y_COORD_21_166_0: value  <=  0;
            Y_COORD_21_166_1: value  <=  0;
            Y_COORD_21_166_2: value  <=  2;
            Y_COORD_21_167_0: value  <=  0;
            Y_COORD_21_167_1: value  <=  0;
            Y_COORD_21_168_0: value  <=  16;
            Y_COORD_21_168_1: value  <=  17;
            Y_COORD_21_169_0: value  <=  4;
            Y_COORD_21_169_1: value  <=  9;
            Y_COORD_21_170_0: value  <=  10;
            Y_COORD_21_170_1: value  <=  11;
            Y_COORD_21_171_0: value  <=  5;
            Y_COORD_21_171_1: value  <=  8;
            Y_COORD_21_172_0: value  <=  0;
            Y_COORD_21_172_1: value  <=  0;
            Y_COORD_21_173_0: value  <=  6;
            Y_COORD_21_173_1: value  <=  6;
            Y_COORD_21_173_2: value  <=  12;
            Y_COORD_21_174_0: value  <=  2;
            Y_COORD_21_174_1: value  <=  4;
            Y_COORD_21_175_0: value  <=  15;
            Y_COORD_21_175_1: value  <=  16;
            Y_COORD_21_176_0: value  <=  0;
            Y_COORD_21_176_1: value  <=  0;
            Y_COORD_21_177_0: value  <=  5;
            Y_COORD_21_177_1: value  <=  5;
            Y_COORD_21_178_0: value  <=  5;
            Y_COORD_21_178_1: value  <=  5;
            Y_COORD_21_179_0: value  <=  6;
            Y_COORD_21_179_1: value  <=  6;
            Y_COORD_21_180_0: value  <=  14;
            Y_COORD_21_180_1: value  <=  14;
            Y_COORD_21_180_2: value  <=  16;
            Y_COORD_21_181_0: value  <=  14;
            Y_COORD_21_181_1: value  <=  14;
            Y_COORD_21_181_2: value  <=  17;
            Y_COORD_21_182_0: value  <=  8;
            Y_COORD_21_182_1: value  <=  12;
            Y_COORD_21_183_0: value  <=  0;
            Y_COORD_21_183_1: value  <=  0;
            Y_COORD_21_183_2: value  <=  4;
            Y_COORD_21_184_0: value  <=  0;
            Y_COORD_21_184_1: value  <=  0;
            Y_COORD_21_184_2: value  <=  4;
            Y_COORD_21_185_0: value  <=  1;
            Y_COORD_21_185_1: value  <=  2;
            Y_COORD_21_186_0: value  <=  9;
            Y_COORD_21_186_1: value  <=  14;
            Y_COORD_21_187_0: value  <=  14;
            Y_COORD_21_187_1: value  <=  15;
            Y_COORD_21_188_0: value  <=  7;
            Y_COORD_21_188_1: value  <=  11;
            Y_COORD_21_189_0: value  <=  7;
            Y_COORD_21_189_1: value  <=  10;
            Y_COORD_21_190_0: value  <=  13;
            Y_COORD_21_190_1: value  <=  14;
            Y_COORD_21_191_0: value  <=  9;
            Y_COORD_21_191_1: value  <=  10;
            Y_COORD_21_192_0: value  <=  1;
            Y_COORD_21_192_1: value  <=  1;
            Y_COORD_21_193_0: value  <=  1;
            Y_COORD_21_193_1: value  <=  8;
            Y_COORD_21_194_0: value  <=  9;
            Y_COORD_21_194_1: value  <=  9;
            Y_COORD_21_195_0: value  <=  7;
            Y_COORD_21_195_1: value  <=  7;
            Y_COORD_21_196_0: value  <=  3;
            Y_COORD_21_196_1: value  <=  3;
            Y_COORD_21_197_0: value  <=  14;
            Y_COORD_21_197_1: value  <=  15;
            Y_COORD_21_198_0: value  <=  11;
            Y_COORD_21_198_1: value  <=  11;
            Y_COORD_21_199_0: value  <=  8;
            Y_COORD_21_199_1: value  <=  8;
            Y_COORD_21_200_0: value  <=  14;
            Y_COORD_21_200_1: value  <=  14;
            Y_COORD_21_201_0: value  <=  8;
            Y_COORD_21_201_1: value  <=  8;
            Y_COORD_21_202_0: value  <=  8;
            Y_COORD_21_202_1: value  <=  8;
            Y_COORD_21_203_0: value  <=  9;
            Y_COORD_21_203_1: value  <=  12;
            Y_COORD_21_204_0: value  <=  14;
            Y_COORD_21_204_1: value  <=  15;
            Y_COORD_21_205_0: value  <=  12;
            Y_COORD_21_205_1: value  <=  13;
            Y_COORD_21_206_0: value  <=  3;
            Y_COORD_21_206_1: value  <=  3;
            Y_COORD_21_207_0: value  <=  4;
            Y_COORD_21_207_1: value  <=  4;
            Y_COORD_21_208_0: value  <=  14;
            Y_COORD_21_208_1: value  <=  15;
            Y_COORD_21_209_0: value  <=  14;
            Y_COORD_21_209_1: value  <=  15;
            Y_COORD_21_210_0: value  <=  15;
            Y_COORD_21_210_1: value  <=  17;
            Y_COORD_21_211_0: value  <=  14;
            Y_COORD_21_211_1: value  <=  17;
            Y_COORD_21_212_0: value  <=  0;
            Y_COORD_21_212_1: value  <=  0;
            Y_COORD_21_212_2: value  <=  3;

            default: value <= 0;

        endcase

    end

endmodule 
