module Height (

input int stage_num,
input int feature_num,
input int rectangle_num,
output real value

);

string name;
assign name = {"HEIGHT_", $sformatf("%d", stage_num),
					"_", $sformatf("%d", feature_num), "_",
					$sformatf("%d", rectangle_num)};

always_comb
    begin

        case (name)

            "HEIGHT_0_0_0": value  <=  4;
            "HEIGHT_0_0_1": value  <=  2;
            "HEIGHT_0_1_0": value  <=  4;
            "HEIGHT_0_1_1": value  <=  4;
            "HEIGHT_0_2_0": value  <=  9;
            "HEIGHT_0_2_1": value  <=  3;
            "HEIGHT_1_0_0": value  <=  6;
            "HEIGHT_1_0_1": value  <=  3;
            "HEIGHT_1_1_0": value  <=  3;
            "HEIGHT_1_1_1": value  <=  3;
            "HEIGHT_1_2_0": value  <=  9;
            "HEIGHT_1_2_1": value  <=  3;
            "HEIGHT_1_3_0": value  <=  8;
            "HEIGHT_1_3_1": value  <=  4;
            "HEIGHT_1_4_0": value  <=  8;
            "HEIGHT_1_4_1": value  <=  4;
            "HEIGHT_1_5_0": value  <=  10;
            "HEIGHT_1_5_1": value  <=  10;
            "HEIGHT_1_6_0": value  <=  12;
            "HEIGHT_1_6_1": value  <=  4;
            "HEIGHT_1_7_0": value  <=  3;
            "HEIGHT_1_7_1": value  <=  3;
            "HEIGHT_1_8_0": value  <=  2;
            "HEIGHT_1_8_1": value  <=  1;
            "HEIGHT_1_9_0": value  <=  2;
            "HEIGHT_1_9_1": value  <=  1;
            "HEIGHT_1_10_0": value  <=  2;
            "HEIGHT_1_10_1": value  <=  1;
            "HEIGHT_1_11_0": value  <=  12;
            "HEIGHT_1_11_1": value  <=  12;
            "HEIGHT_1_12_0": value  <=  12;
            "HEIGHT_1_12_1": value  <=  6;
            "HEIGHT_1_12_2": value  <=  6;
            "HEIGHT_1_13_0": value  <=  8;
            "HEIGHT_1_13_1": value  <=  8;
            "HEIGHT_1_14_0": value  <=  2;
            "HEIGHT_1_14_1": value  <=  1;
            "HEIGHT_1_15_0": value  <=  3;
            "HEIGHT_1_15_1": value  <=  1;
            "HEIGHT_2_0_0": value  <=  9;
            "HEIGHT_2_0_1": value  <=  3;
            "HEIGHT_2_1_0": value  <=  14;
            "HEIGHT_2_1_1": value  <=  7;
            "HEIGHT_2_2_0": value  <=  12;
            "HEIGHT_2_2_1": value  <=  4;
            "HEIGHT_2_3_0": value  <=  5;
            "HEIGHT_2_3_1": value  <=  5;
            "HEIGHT_2_4_0": value  <=  8;
            "HEIGHT_2_4_1": value  <=  4;
            "HEIGHT_2_5_0": value  <=  9;
            "HEIGHT_2_5_1": value  <=  3;
            "HEIGHT_2_6_0": value  <=  8;
            "HEIGHT_2_6_1": value  <=  4;
            "HEIGHT_2_7_0": value  <=  6;
            "HEIGHT_2_7_1": value  <=  2;
            "HEIGHT_2_8_0": value  <=  17;
            "HEIGHT_2_8_1": value  <=  17;
            "HEIGHT_2_9_0": value  <=  4;
            "HEIGHT_2_9_1": value  <=  4;
            "HEIGHT_2_10_0": value  <=  4;
            "HEIGHT_2_10_1": value  <=  4;
            "HEIGHT_2_11_0": value  <=  16;
            "HEIGHT_2_11_1": value  <=  16;
            "HEIGHT_2_12_0": value  <=  8;
            "HEIGHT_2_12_1": value  <=  4;
            "HEIGHT_2_12_2": value  <=  4;
            "HEIGHT_2_13_0": value  <=  4;
            "HEIGHT_2_13_1": value  <=  2;
            "HEIGHT_2_13_2": value  <=  2;
            "HEIGHT_2_14_0": value  <=  8;
            "HEIGHT_2_14_1": value  <=  4;
            "HEIGHT_2_14_2": value  <=  4;
            "HEIGHT_2_15_0": value  <=  10;
            "HEIGHT_2_15_1": value  <=  5;
            "HEIGHT_2_15_2": value  <=  5;
            "HEIGHT_2_16_0": value  <=  16;
            "HEIGHT_2_16_1": value  <=  16;
            "HEIGHT_2_17_0": value  <=  2;
            "HEIGHT_2_17_1": value  <=  1;
            "HEIGHT_2_18_0": value  <=  3;
            "HEIGHT_2_18_1": value  <=  1;
            "HEIGHT_2_19_0": value  <=  3;
            "HEIGHT_2_19_1": value  <=  1;
            "HEIGHT_2_20_0": value  <=  6;
            "HEIGHT_2_20_1": value  <=  2;
            "HEIGHT_3_0_0": value  <=  4;
            "HEIGHT_3_0_1": value  <=  2;
            "HEIGHT_3_1_0": value  <=  16;
            "HEIGHT_3_1_1": value  <=  8;
            "HEIGHT_3_2_0": value  <=  8;
            "HEIGHT_3_2_1": value  <=  4;
            "HEIGHT_3_3_0": value  <=  2;
            "HEIGHT_3_3_1": value  <=  2;
            "HEIGHT_3_4_0": value  <=  12;
            "HEIGHT_3_4_1": value  <=  4;
            "HEIGHT_3_5_0": value  <=  6;
            "HEIGHT_3_5_1": value  <=  3;
            "HEIGHT_3_5_2": value  <=  3;
            "HEIGHT_3_6_0": value  <=  19;
            "HEIGHT_3_6_1": value  <=  19;
            "HEIGHT_3_7_0": value  <=  4;
            "HEIGHT_3_7_1": value  <=  4;
            "HEIGHT_3_8_0": value  <=  3;
            "HEIGHT_3_8_1": value  <=  3;
            "HEIGHT_3_9_0": value  <=  4;
            "HEIGHT_3_9_1": value  <=  2;
            "HEIGHT_3_9_2": value  <=  2;
            "HEIGHT_3_10_0": value  <=  10;
            "HEIGHT_3_10_1": value  <=  10;
            "HEIGHT_3_11_0": value  <=  15;
            "HEIGHT_3_11_1": value  <=  5;
            "HEIGHT_3_12_0": value  <=  6;
            "HEIGHT_3_12_1": value  <=  2;
            "HEIGHT_3_13_0": value  <=  10;
            "HEIGHT_3_13_1": value  <=  5;
            "HEIGHT_3_13_2": value  <=  5;
            "HEIGHT_3_14_0": value  <=  4;
            "HEIGHT_3_14_1": value  <=  4;
            "HEIGHT_3_15_0": value  <=  2;
            "HEIGHT_3_15_1": value  <=  1;
            "HEIGHT_3_16_0": value  <=  2;
            "HEIGHT_3_16_1": value  <=  1;
            "HEIGHT_3_17_0": value  <=  3;
            "HEIGHT_3_17_1": value  <=  1;
            "HEIGHT_3_18_0": value  <=  4;
            "HEIGHT_3_18_1": value  <=  2;
            "HEIGHT_3_18_2": value  <=  2;
            "HEIGHT_3_19_0": value  <=  2;
            "HEIGHT_3_19_1": value  <=  1;
            "HEIGHT_3_20_0": value  <=  3;
            "HEIGHT_3_20_1": value  <=  1;
            "HEIGHT_3_21_0": value  <=  2;
            "HEIGHT_3_21_1": value  <=  1;
            "HEIGHT_3_22_0": value  <=  3;
            "HEIGHT_3_22_1": value  <=  1;
            "HEIGHT_3_23_0": value  <=  2;
            "HEIGHT_3_23_1": value  <=  1;
            "HEIGHT_3_24_0": value  <=  6;
            "HEIGHT_3_24_1": value  <=  2;
            "HEIGHT_3_25_0": value  <=  2;
            "HEIGHT_3_25_1": value  <=  2;
            "HEIGHT_3_26_0": value  <=  9;
            "HEIGHT_3_26_1": value  <=  3;
            "HEIGHT_3_27_0": value  <=  2;
            "HEIGHT_3_27_1": value  <=  2;
            "HEIGHT_3_28_0": value  <=  2;
            "HEIGHT_3_28_1": value  <=  1;
            "HEIGHT_3_29_0": value  <=  4;
            "HEIGHT_3_29_1": value  <=  4;
            "HEIGHT_3_30_0": value  <=  2;
            "HEIGHT_3_30_1": value  <=  2;
            "HEIGHT_3_31_0": value  <=  3;
            "HEIGHT_3_31_1": value  <=  3;
            "HEIGHT_3_32_0": value  <=  2;
            "HEIGHT_3_32_1": value  <=  1;
            "HEIGHT_3_33_0": value  <=  2;
            "HEIGHT_3_33_1": value  <=  2;
            "HEIGHT_3_34_0": value  <=  4;
            "HEIGHT_3_34_1": value  <=  2;
            "HEIGHT_3_35_0": value  <=  4;
            "HEIGHT_3_35_1": value  <=  2;
            "HEIGHT_3_35_2": value  <=  2;
            "HEIGHT_3_36_0": value  <=  3;
            "HEIGHT_3_36_1": value  <=  1;
            "HEIGHT_3_37_0": value  <=  6;
            "HEIGHT_3_37_1": value  <=  6;
            "HEIGHT_3_38_0": value  <=  6;
            "HEIGHT_3_38_1": value  <=  6;
            "HEIGHT_4_0_0": value  <=  9;
            "HEIGHT_4_0_1": value  <=  3;
            "HEIGHT_4_1_0": value  <=  6;
            "HEIGHT_4_1_1": value  <=  3;
            "HEIGHT_4_2_0": value  <=  8;
            "HEIGHT_4_2_1": value  <=  4;
            "HEIGHT_4_3_0": value  <=  9;
            "HEIGHT_4_3_1": value  <=  9;
            "HEIGHT_4_4_0": value  <=  1;
            "HEIGHT_4_4_1": value  <=  1;
            "HEIGHT_4_5_0": value  <=  1;
            "HEIGHT_4_5_1": value  <=  1;
            "HEIGHT_4_6_0": value  <=  6;
            "HEIGHT_4_6_1": value  <=  3;
            "HEIGHT_4_7_0": value  <=  1;
            "HEIGHT_4_7_1": value  <=  1;
            "HEIGHT_4_8_0": value  <=  6;
            "HEIGHT_4_8_1": value  <=  2;
            "HEIGHT_4_9_0": value  <=  6;
            "HEIGHT_4_9_1": value  <=  2;
            "HEIGHT_4_10_0": value  <=  2;
            "HEIGHT_4_10_1": value  <=  2;
            "HEIGHT_4_11_0": value  <=  1;
            "HEIGHT_4_11_1": value  <=  1;
            "HEIGHT_4_12_0": value  <=  14;
            "HEIGHT_4_12_1": value  <=  14;
            "HEIGHT_4_13_0": value  <=  4;
            "HEIGHT_4_13_1": value  <=  2;
            "HEIGHT_4_13_2": value  <=  2;
            "HEIGHT_4_14_0": value  <=  14;
            "HEIGHT_4_14_1": value  <=  7;
            "HEIGHT_4_15_0": value  <=  4;
            "HEIGHT_4_15_1": value  <=  2;
            "HEIGHT_4_16_0": value  <=  4;
            "HEIGHT_4_16_1": value  <=  4;
            "HEIGHT_4_17_0": value  <=  2;
            "HEIGHT_4_17_1": value  <=  2;
            "HEIGHT_4_18_0": value  <=  2;
            "HEIGHT_4_18_1": value  <=  2;
            "HEIGHT_4_19_0": value  <=  6;
            "HEIGHT_4_19_1": value  <=  2;
            "HEIGHT_4_20_0": value  <=  6;
            "HEIGHT_4_20_1": value  <=  2;
            "HEIGHT_4_21_0": value  <=  12;
            "HEIGHT_4_21_1": value  <=  4;
            "HEIGHT_4_22_0": value  <=  2;
            "HEIGHT_4_22_1": value  <=  2;
            "HEIGHT_4_23_0": value  <=  2;
            "HEIGHT_4_23_1": value  <=  2;
            "HEIGHT_4_24_0": value  <=  3;
            "HEIGHT_4_24_1": value  <=  1;
            "HEIGHT_4_25_0": value  <=  2;
            "HEIGHT_4_25_1": value  <=  2;
            "HEIGHT_4_26_0": value  <=  5;
            "HEIGHT_4_26_1": value  <=  5;
            "HEIGHT_4_27_0": value  <=  4;
            "HEIGHT_4_27_1": value  <=  2;
            "HEIGHT_4_27_2": value  <=  2;
            "HEIGHT_4_28_0": value  <=  3;
            "HEIGHT_4_28_1": value  <=  1;
            "HEIGHT_4_29_0": value  <=  3;
            "HEIGHT_4_29_1": value  <=  1;
            "HEIGHT_4_30_0": value  <=  12;
            "HEIGHT_4_30_1": value  <=  6;
            "HEIGHT_4_30_2": value  <=  6;
            "HEIGHT_4_31_0": value  <=  12;
            "HEIGHT_4_31_1": value  <=  4;
            "HEIGHT_4_32_0": value  <=  14;
            "HEIGHT_4_32_1": value  <=  7;
            "HEIGHT_4_32_2": value  <=  7;
            "HEIGHT_5_0_0": value  <=  2;
            "HEIGHT_5_0_1": value  <=  2;
            "HEIGHT_5_1_0": value  <=  4;
            "HEIGHT_5_1_1": value  <=  2;
            "HEIGHT_5_2_0": value  <=  8;
            "HEIGHT_5_2_1": value  <=  4;
            "HEIGHT_5_3_0": value  <=  4;
            "HEIGHT_5_3_1": value  <=  2;
            "HEIGHT_5_4_0": value  <=  2;
            "HEIGHT_5_4_1": value  <=  1;
            "HEIGHT_5_5_0": value  <=  2;
            "HEIGHT_5_5_1": value  <=  2;
            "HEIGHT_5_6_0": value  <=  10;
            "HEIGHT_5_6_1": value  <=  5;
            "HEIGHT_5_6_2": value  <=  5;
            "HEIGHT_5_7_0": value  <=  15;
            "HEIGHT_5_7_1": value  <=  5;
            "HEIGHT_5_8_0": value  <=  6;
            "HEIGHT_5_8_1": value  <=  3;
            "HEIGHT_5_8_2": value  <=  3;
            "HEIGHT_5_9_0": value  <=  2;
            "HEIGHT_5_9_1": value  <=  1;
            "HEIGHT_5_10_0": value  <=  6;
            "HEIGHT_5_10_1": value  <=  3;
            "HEIGHT_5_11_0": value  <=  3;
            "HEIGHT_5_11_1": value  <=  3;
            "HEIGHT_5_12_0": value  <=  6;
            "HEIGHT_5_12_1": value  <=  3;
            "HEIGHT_5_12_2": value  <=  3;
            "HEIGHT_5_13_0": value  <=  4;
            "HEIGHT_5_13_1": value  <=  2;
            "HEIGHT_5_14_0": value  <=  8;
            "HEIGHT_5_14_1": value  <=  4;
            "HEIGHT_5_14_2": value  <=  4;
            "HEIGHT_5_15_0": value  <=  2;
            "HEIGHT_5_15_1": value  <=  1;
            "HEIGHT_5_16_0": value  <=  2;
            "HEIGHT_5_16_1": value  <=  2;
            "HEIGHT_5_17_0": value  <=  8;
            "HEIGHT_5_17_1": value  <=  4;
            "HEIGHT_5_18_0": value  <=  3;
            "HEIGHT_5_18_1": value  <=  1;
            "HEIGHT_5_19_0": value  <=  8;
            "HEIGHT_5_19_1": value  <=  4;
            "HEIGHT_5_19_2": value  <=  4;
            "HEIGHT_5_20_0": value  <=  6;
            "HEIGHT_5_20_1": value  <=  3;
            "HEIGHT_5_21_0": value  <=  3;
            "HEIGHT_5_21_1": value  <=  1;
            "HEIGHT_5_22_0": value  <=  6;
            "HEIGHT_5_22_1": value  <=  6;
            "HEIGHT_5_23_0": value  <=  3;
            "HEIGHT_5_23_1": value  <=  1;
            "HEIGHT_5_24_0": value  <=  3;
            "HEIGHT_5_24_1": value  <=  1;
            "HEIGHT_5_25_0": value  <=  12;
            "HEIGHT_5_25_1": value  <=  6;
            "HEIGHT_5_25_2": value  <=  6;
            "HEIGHT_5_26_0": value  <=  3;
            "HEIGHT_5_26_1": value  <=  3;
            "HEIGHT_5_27_0": value  <=  10;
            "HEIGHT_5_27_1": value  <=  5;
            "HEIGHT_5_28_0": value  <=  12;
            "HEIGHT_5_28_1": value  <=  12;
            "HEIGHT_5_29_0": value  <=  3;
            "HEIGHT_5_29_1": value  <=  1;
            "HEIGHT_5_30_0": value  <=  3;
            "HEIGHT_5_30_1": value  <=  1;
            "HEIGHT_5_31_0": value  <=  3;
            "HEIGHT_5_31_1": value  <=  1;
            "HEIGHT_5_32_0": value  <=  3;
            "HEIGHT_5_32_1": value  <=  1;
            "HEIGHT_5_33_0": value  <=  3;
            "HEIGHT_5_33_1": value  <=  1;
            "HEIGHT_5_34_0": value  <=  3;
            "HEIGHT_5_34_1": value  <=  1;
            "HEIGHT_5_35_0": value  <=  12;
            "HEIGHT_5_35_1": value  <=  6;
            "HEIGHT_5_35_2": value  <=  6;
            "HEIGHT_5_36_0": value  <=  6;
            "HEIGHT_5_36_1": value  <=  6;
            "HEIGHT_5_37_0": value  <=  2;
            "HEIGHT_5_37_1": value  <=  1;
            "HEIGHT_5_38_0": value  <=  4;
            "HEIGHT_5_38_1": value  <=  4;
            "HEIGHT_5_39_0": value  <=  8;
            "HEIGHT_5_39_1": value  <=  4;
            "HEIGHT_5_40_0": value  <=  6;
            "HEIGHT_5_40_1": value  <=  6;
            "HEIGHT_5_41_0": value  <=  3;
            "HEIGHT_5_41_1": value  <=  3;
            "HEIGHT_5_42_0": value  <=  1;
            "HEIGHT_5_42_1": value  <=  1;
            "HEIGHT_5_43_0": value  <=  3;
            "HEIGHT_5_43_1": value  <=  1;
            "HEIGHT_6_0_0": value  <=  9;
            "HEIGHT_6_0_1": value  <=  3;
            "HEIGHT_6_1_0": value  <=  1;
            "HEIGHT_6_1_1": value  <=  1;
            "HEIGHT_6_2_0": value  <=  8;
            "HEIGHT_6_2_1": value  <=  4;
            "HEIGHT_6_3_0": value  <=  6;
            "HEIGHT_6_3_1": value  <=  3;
            "HEIGHT_6_4_0": value  <=  15;
            "HEIGHT_6_4_1": value  <=  5;
            "HEIGHT_6_5_0": value  <=  9;
            "HEIGHT_6_5_1": value  <=  3;
            "HEIGHT_6_6_0": value  <=  14;
            "HEIGHT_6_6_1": value  <=  7;
            "HEIGHT_6_7_0": value  <=  6;
            "HEIGHT_6_7_1": value  <=  2;
            "HEIGHT_6_8_0": value  <=  4;
            "HEIGHT_6_8_1": value  <=  4;
            "HEIGHT_6_9_0": value  <=  10;
            "HEIGHT_6_9_1": value  <=  5;
            "HEIGHT_6_10_0": value  <=  6;
            "HEIGHT_6_10_1": value  <=  2;
            "HEIGHT_6_11_0": value  <=  10;
            "HEIGHT_6_11_1": value  <=  10;
            "HEIGHT_6_12_0": value  <=  10;
            "HEIGHT_6_12_1": value  <=  5;
            "HEIGHT_6_12_2": value  <=  5;
            "HEIGHT_6_13_0": value  <=  12;
            "HEIGHT_6_13_1": value  <=  6;
            "HEIGHT_6_13_2": value  <=  6;
            "HEIGHT_6_14_0": value  <=  9;
            "HEIGHT_6_14_1": value  <=  9;
            "HEIGHT_6_15_0": value  <=  5;
            "HEIGHT_6_15_1": value  <=  5;
            "HEIGHT_6_16_0": value  <=  5;
            "HEIGHT_6_16_1": value  <=  5;
            "HEIGHT_6_17_0": value  <=  3;
            "HEIGHT_6_17_1": value  <=  1;
            "HEIGHT_6_18_0": value  <=  2;
            "HEIGHT_6_18_1": value  <=  2;
            "HEIGHT_6_19_0": value  <=  3;
            "HEIGHT_6_19_1": value  <=  1;
            "HEIGHT_6_20_0": value  <=  6;
            "HEIGHT_6_20_1": value  <=  3;
            "HEIGHT_6_21_0": value  <=  9;
            "HEIGHT_6_21_1": value  <=  3;
            "HEIGHT_6_22_0": value  <=  2;
            "HEIGHT_6_22_1": value  <=  1;
            "HEIGHT_6_23_0": value  <=  5;
            "HEIGHT_6_23_1": value  <=  5;
            "HEIGHT_6_24_0": value  <=  7;
            "HEIGHT_6_24_1": value  <=  7;
            "HEIGHT_6_25_0": value  <=  9;
            "HEIGHT_6_25_1": value  <=  3;
            "HEIGHT_6_26_0": value  <=  8;
            "HEIGHT_6_26_1": value  <=  4;
            "HEIGHT_6_26_2": value  <=  4;
            "HEIGHT_6_27_0": value  <=  6;
            "HEIGHT_6_27_1": value  <=  2;
            "HEIGHT_6_28_0": value  <=  6;
            "HEIGHT_6_28_1": value  <=  2;
            "HEIGHT_6_29_0": value  <=  4;
            "HEIGHT_6_29_1": value  <=  2;
            "HEIGHT_6_30_0": value  <=  3;
            "HEIGHT_6_30_1": value  <=  1;
            "HEIGHT_6_31_0": value  <=  8;
            "HEIGHT_6_31_1": value  <=  4;
            "HEIGHT_6_32_0": value  <=  4;
            "HEIGHT_6_32_1": value  <=  4;
            "HEIGHT_6_33_0": value  <=  1;
            "HEIGHT_6_33_1": value  <=  1;
            "HEIGHT_6_34_0": value  <=  3;
            "HEIGHT_6_34_1": value  <=  1;
            "HEIGHT_6_35_0": value  <=  6;
            "HEIGHT_6_35_1": value  <=  3;
            "HEIGHT_6_35_2": value  <=  3;
            "HEIGHT_6_36_0": value  <=  5;
            "HEIGHT_6_36_1": value  <=  5;
            "HEIGHT_6_37_0": value  <=  3;
            "HEIGHT_6_37_1": value  <=  1;
            "HEIGHT_6_38_0": value  <=  2;
            "HEIGHT_6_38_1": value  <=  1;
            "HEIGHT_6_39_0": value  <=  3;
            "HEIGHT_6_39_1": value  <=  1;
            "HEIGHT_6_40_0": value  <=  4;
            "HEIGHT_6_40_1": value  <=  4;
            "HEIGHT_6_41_0": value  <=  8;
            "HEIGHT_6_41_1": value  <=  8;
            "HEIGHT_6_42_0": value  <=  2;
            "HEIGHT_6_42_1": value  <=  2;
            "HEIGHT_6_43_0": value  <=  4;
            "HEIGHT_6_43_1": value  <=  2;
            "HEIGHT_6_43_2": value  <=  2;
            "HEIGHT_6_44_0": value  <=  6;
            "HEIGHT_6_44_1": value  <=  2;
            "HEIGHT_6_45_0": value  <=  4;
            "HEIGHT_6_45_1": value  <=  2;
            "HEIGHT_6_46_0": value  <=  4;
            "HEIGHT_6_46_1": value  <=  2;
            "HEIGHT_6_47_0": value  <=  8;
            "HEIGHT_6_47_1": value  <=  4;
            "HEIGHT_6_47_2": value  <=  4;
            "HEIGHT_6_48_0": value  <=  3;
            "HEIGHT_6_48_1": value  <=  1;
            "HEIGHT_6_49_0": value  <=  4;
            "HEIGHT_6_49_1": value  <=  2;
            "HEIGHT_7_0_0": value  <=  1;
            "HEIGHT_7_0_1": value  <=  1;
            "HEIGHT_7_1_0": value  <=  6;
            "HEIGHT_7_1_1": value  <=  3;
            "HEIGHT_7_1_2": value  <=  3;
            "HEIGHT_7_2_0": value  <=  6;
            "HEIGHT_7_2_1": value  <=  2;
            "HEIGHT_7_3_0": value  <=  14;
            "HEIGHT_7_3_1": value  <=  7;
            "HEIGHT_7_3_2": value  <=  7;
            "HEIGHT_7_4_0": value  <=  15;
            "HEIGHT_7_4_1": value  <=  5;
            "HEIGHT_7_5_0": value  <=  8;
            "HEIGHT_7_5_1": value  <=  4;
            "HEIGHT_7_5_2": value  <=  4;
            "HEIGHT_7_6_0": value  <=  8;
            "HEIGHT_7_6_1": value  <=  4;
            "HEIGHT_7_6_2": value  <=  4;
            "HEIGHT_7_7_0": value  <=  7;
            "HEIGHT_7_7_1": value  <=  7;
            "HEIGHT_7_8_0": value  <=  14;
            "HEIGHT_7_8_1": value  <=  7;
            "HEIGHT_7_8_2": value  <=  7;
            "HEIGHT_7_9_0": value  <=  6;
            "HEIGHT_7_9_1": value  <=  2;
            "HEIGHT_7_10_0": value  <=  3;
            "HEIGHT_7_10_1": value  <=  1;
            "HEIGHT_7_11_0": value  <=  6;
            "HEIGHT_7_11_1": value  <=  2;
            "HEIGHT_7_12_0": value  <=  6;
            "HEIGHT_7_12_1": value  <=  2;
            "HEIGHT_7_13_0": value  <=  6;
            "HEIGHT_7_13_1": value  <=  2;
            "HEIGHT_7_14_0": value  <=  7;
            "HEIGHT_7_14_1": value  <=  7;
            "HEIGHT_7_15_0": value  <=  14;
            "HEIGHT_7_15_1": value  <=  7;
            "HEIGHT_7_16_0": value  <=  10;
            "HEIGHT_7_16_1": value  <=  5;
            "HEIGHT_7_17_0": value  <=  2;
            "HEIGHT_7_17_1": value  <=  1;
            "HEIGHT_7_18_0": value  <=  4;
            "HEIGHT_7_18_1": value  <=  2;
            "HEIGHT_7_18_2": value  <=  2;
            "HEIGHT_7_19_0": value  <=  4;
            "HEIGHT_7_19_1": value  <=  2;
            "HEIGHT_7_19_2": value  <=  2;
            "HEIGHT_7_20_0": value  <=  9;
            "HEIGHT_7_20_1": value  <=  3;
            "HEIGHT_7_21_0": value  <=  6;
            "HEIGHT_7_21_1": value  <=  3;
            "HEIGHT_7_22_0": value  <=  1;
            "HEIGHT_7_22_1": value  <=  1;
            "HEIGHT_7_23_0": value  <=  5;
            "HEIGHT_7_23_1": value  <=  5;
            "HEIGHT_7_24_0": value  <=  4;
            "HEIGHT_7_24_1": value  <=  2;
            "HEIGHT_7_25_0": value  <=  6;
            "HEIGHT_7_25_1": value  <=  2;
            "HEIGHT_7_26_0": value  <=  2;
            "HEIGHT_7_26_1": value  <=  2;
            "HEIGHT_7_27_0": value  <=  2;
            "HEIGHT_7_27_1": value  <=  2;
            "HEIGHT_7_28_0": value  <=  2;
            "HEIGHT_7_28_1": value  <=  2;
            "HEIGHT_7_29_0": value  <=  2;
            "HEIGHT_7_29_1": value  <=  1;
            "HEIGHT_7_30_0": value  <=  3;
            "HEIGHT_7_30_1": value  <=  1;
            "HEIGHT_7_31_0": value  <=  4;
            "HEIGHT_7_31_1": value  <=  4;
            "HEIGHT_7_32_0": value  <=  3;
            "HEIGHT_7_32_1": value  <=  1;
            "HEIGHT_7_33_0": value  <=  6;
            "HEIGHT_7_33_1": value  <=  3;
            "HEIGHT_7_33_2": value  <=  3;
            "HEIGHT_7_34_0": value  <=  3;
            "HEIGHT_7_34_1": value  <=  1;
            "HEIGHT_7_35_0": value  <=  3;
            "HEIGHT_7_35_1": value  <=  1;
            "HEIGHT_7_36_0": value  <=  8;
            "HEIGHT_7_36_1": value  <=  8;
            "HEIGHT_7_37_0": value  <=  6;
            "HEIGHT_7_37_1": value  <=  6;
            "HEIGHT_7_38_0": value  <=  8;
            "HEIGHT_7_38_1": value  <=  8;
            "HEIGHT_7_39_0": value  <=  13;
            "HEIGHT_7_39_1": value  <=  13;
            "HEIGHT_7_40_0": value  <=  6;
            "HEIGHT_7_40_1": value  <=  3;
            "HEIGHT_7_41_0": value  <=  13;
            "HEIGHT_7_41_1": value  <=  13;
            "HEIGHT_7_42_0": value  <=  4;
            "HEIGHT_7_42_1": value  <=  2;
            "HEIGHT_7_42_2": value  <=  2;
            "HEIGHT_7_43_0": value  <=  13;
            "HEIGHT_7_43_1": value  <=  13;
            "HEIGHT_7_44_0": value  <=  13;
            "HEIGHT_7_44_1": value  <=  13;
            "HEIGHT_7_45_0": value  <=  1;
            "HEIGHT_7_45_1": value  <=  1;
            "HEIGHT_7_46_0": value  <=  1;
            "HEIGHT_7_46_1": value  <=  1;
            "HEIGHT_7_47_0": value  <=  4;
            "HEIGHT_7_47_1": value  <=  2;
            "HEIGHT_7_47_2": value  <=  2;
            "HEIGHT_7_48_0": value  <=  3;
            "HEIGHT_7_48_1": value  <=  3;
            "HEIGHT_7_49_0": value  <=  2;
            "HEIGHT_7_49_1": value  <=  2;
            "HEIGHT_7_50_0": value  <=  5;
            "HEIGHT_7_50_1": value  <=  5;
            "HEIGHT_8_0_0": value  <=  6;
            "HEIGHT_8_0_1": value  <=  2;
            "HEIGHT_8_1_0": value  <=  12;
            "HEIGHT_8_1_1": value  <=  6;
            "HEIGHT_8_2_0": value  <=  8;
            "HEIGHT_8_2_1": value  <=  4;
            "HEIGHT_8_3_0": value  <=  5;
            "HEIGHT_8_3_1": value  <=  5;
            "HEIGHT_8_4_0": value  <=  3;
            "HEIGHT_8_4_1": value  <=  1;
            "HEIGHT_8_5_0": value  <=  8;
            "HEIGHT_8_5_1": value  <=  4;
            "HEIGHT_8_6_0": value  <=  5;
            "HEIGHT_8_6_1": value  <=  5;
            "HEIGHT_8_7_0": value  <=  4;
            "HEIGHT_8_7_1": value  <=  2;
            "HEIGHT_8_8_0": value  <=  1;
            "HEIGHT_8_8_1": value  <=  1;
            "HEIGHT_8_9_0": value  <=  1;
            "HEIGHT_8_9_1": value  <=  1;
            "HEIGHT_8_10_0": value  <=  3;
            "HEIGHT_8_10_1": value  <=  1;
            "HEIGHT_8_11_0": value  <=  6;
            "HEIGHT_8_11_1": value  <=  3;
            "HEIGHT_8_12_0": value  <=  6;
            "HEIGHT_8_12_1": value  <=  3;
            "HEIGHT_8_13_0": value  <=  6;
            "HEIGHT_8_13_1": value  <=  2;
            "HEIGHT_8_14_0": value  <=  3;
            "HEIGHT_8_14_1": value  <=  1;
            "HEIGHT_8_15_0": value  <=  5;
            "HEIGHT_8_15_1": value  <=  5;
            "HEIGHT_8_16_0": value  <=  9;
            "HEIGHT_8_16_1": value  <=  9;
            "HEIGHT_8_17_0": value  <=  1;
            "HEIGHT_8_17_1": value  <=  1;
            "HEIGHT_8_18_0": value  <=  4;
            "HEIGHT_8_18_1": value  <=  2;
            "HEIGHT_8_19_0": value  <=  2;
            "HEIGHT_8_19_1": value  <=  1;
            "HEIGHT_8_20_0": value  <=  2;
            "HEIGHT_8_20_1": value  <=  1;
            "HEIGHT_8_21_0": value  <=  6;
            "HEIGHT_8_21_1": value  <=  2;
            "HEIGHT_8_22_0": value  <=  2;
            "HEIGHT_8_22_1": value  <=  2;
            "HEIGHT_8_23_0": value  <=  2;
            "HEIGHT_8_23_1": value  <=  1;
            "HEIGHT_8_23_2": value  <=  1;
            "HEIGHT_8_24_0": value  <=  6;
            "HEIGHT_8_24_1": value  <=  3;
            "HEIGHT_8_25_0": value  <=  4;
            "HEIGHT_8_25_1": value  <=  2;
            "HEIGHT_8_25_2": value  <=  2;
            "HEIGHT_8_26_0": value  <=  5;
            "HEIGHT_8_26_1": value  <=  5;
            "HEIGHT_8_27_0": value  <=  2;
            "HEIGHT_8_27_1": value  <=  1;
            "HEIGHT_8_28_0": value  <=  2;
            "HEIGHT_8_28_1": value  <=  1;
            "HEIGHT_8_28_2": value  <=  1;
            "HEIGHT_8_29_0": value  <=  2;
            "HEIGHT_8_29_1": value  <=  1;
            "HEIGHT_8_29_2": value  <=  1;
            "HEIGHT_8_30_0": value  <=  3;
            "HEIGHT_8_30_1": value  <=  1;
            "HEIGHT_8_31_0": value  <=  6;
            "HEIGHT_8_31_1": value  <=  3;
            "HEIGHT_8_31_2": value  <=  3;
            "HEIGHT_8_32_0": value  <=  3;
            "HEIGHT_8_32_1": value  <=  1;
            "HEIGHT_8_33_0": value  <=  6;
            "HEIGHT_8_33_1": value  <=  2;
            "HEIGHT_8_34_0": value  <=  6;
            "HEIGHT_8_34_1": value  <=  2;
            "HEIGHT_8_35_0": value  <=  12;
            "HEIGHT_8_35_1": value  <=  6;
            "HEIGHT_8_35_2": value  <=  6;
            "HEIGHT_8_36_0": value  <=  3;
            "HEIGHT_8_36_1": value  <=  1;
            "HEIGHT_8_37_0": value  <=  3;
            "HEIGHT_8_37_1": value  <=  3;
            "HEIGHT_8_38_0": value  <=  3;
            "HEIGHT_8_38_1": value  <=  1;
            "HEIGHT_8_39_0": value  <=  3;
            "HEIGHT_8_39_1": value  <=  3;
            "HEIGHT_8_40_0": value  <=  10;
            "HEIGHT_8_40_1": value  <=  5;
            "HEIGHT_8_40_2": value  <=  5;
            "HEIGHT_8_41_0": value  <=  2;
            "HEIGHT_8_41_1": value  <=  2;
            "HEIGHT_8_42_0": value  <=  3;
            "HEIGHT_8_42_1": value  <=  3;
            "HEIGHT_8_43_0": value  <=  3;
            "HEIGHT_8_43_1": value  <=  1;
            "HEIGHT_8_44_0": value  <=  4;
            "HEIGHT_8_44_1": value  <=  4;
            "HEIGHT_8_45_0": value  <=  12;
            "HEIGHT_8_45_1": value  <=  6;
            "HEIGHT_8_46_0": value  <=  12;
            "HEIGHT_8_46_1": value  <=  6;
            "HEIGHT_8_46_2": value  <=  6;
            "HEIGHT_8_47_0": value  <=  3;
            "HEIGHT_8_47_1": value  <=  1;
            "HEIGHT_8_48_0": value  <=  3;
            "HEIGHT_8_48_1": value  <=  1;
            "HEIGHT_8_49_0": value  <=  2;
            "HEIGHT_8_49_1": value  <=  1;
            "HEIGHT_8_49_2": value  <=  1;
            "HEIGHT_8_50_0": value  <=  10;
            "HEIGHT_8_50_1": value  <=  10;
            "HEIGHT_8_51_0": value  <=  5;
            "HEIGHT_8_51_1": value  <=  5;
            "HEIGHT_8_52_0": value  <=  2;
            "HEIGHT_8_52_1": value  <=  2;
            "HEIGHT_8_53_0": value  <=  10;
            "HEIGHT_8_53_1": value  <=  5;
            "HEIGHT_8_54_0": value  <=  3;
            "HEIGHT_8_54_1": value  <=  3;
            "HEIGHT_8_55_0": value  <=  6;
            "HEIGHT_8_55_1": value  <=  2;
            "HEIGHT_9_0_0": value  <=  6;
            "HEIGHT_9_0_1": value  <=  3;
            "HEIGHT_9_1_0": value  <=  2;
            "HEIGHT_9_1_1": value  <=  2;
            "HEIGHT_9_2_0": value  <=  10;
            "HEIGHT_9_2_1": value  <=  5;
            "HEIGHT_9_3_0": value  <=  16;
            "HEIGHT_9_3_1": value  <=  8;
            "HEIGHT_9_4_0": value  <=  4;
            "HEIGHT_9_4_1": value  <=  2;
            "HEIGHT_9_5_0": value  <=  9;
            "HEIGHT_9_5_1": value  <=  9;
            "HEIGHT_9_6_0": value  <=  2;
            "HEIGHT_9_6_1": value  <=  1;
            "HEIGHT_9_7_0": value  <=  9;
            "HEIGHT_9_7_1": value  <=  3;
            "HEIGHT_9_8_0": value  <=  3;
            "HEIGHT_9_8_1": value  <=  1;
            "HEIGHT_9_9_0": value  <=  6;
            "HEIGHT_9_9_1": value  <=  3;
            "HEIGHT_9_9_2": value  <=  3;
            "HEIGHT_9_10_0": value  <=  10;
            "HEIGHT_9_10_1": value  <=  5;
            "HEIGHT_9_10_2": value  <=  5;
            "HEIGHT_9_11_0": value  <=  4;
            "HEIGHT_9_11_1": value  <=  2;
            "HEIGHT_9_12_0": value  <=  4;
            "HEIGHT_9_12_1": value  <=  2;
            "HEIGHT_9_13_0": value  <=  3;
            "HEIGHT_9_13_1": value  <=  3;
            "HEIGHT_9_14_0": value  <=  8;
            "HEIGHT_9_14_1": value  <=  4;
            "HEIGHT_9_15_0": value  <=  6;
            "HEIGHT_9_15_1": value  <=  3;
            "HEIGHT_9_16_0": value  <=  6;
            "HEIGHT_9_16_1": value  <=  3;
            "HEIGHT_9_16_2": value  <=  3;
            "HEIGHT_9_17_0": value  <=  12;
            "HEIGHT_9_17_1": value  <=  6;
            "HEIGHT_9_17_2": value  <=  6;
            "HEIGHT_9_18_0": value  <=  2;
            "HEIGHT_9_18_1": value  <=  1;
            "HEIGHT_9_19_0": value  <=  3;
            "HEIGHT_9_19_1": value  <=  1;
            "HEIGHT_9_20_0": value  <=  2;
            "HEIGHT_9_20_1": value  <=  1;
            "HEIGHT_9_21_0": value  <=  3;
            "HEIGHT_9_21_1": value  <=  1;
            "HEIGHT_9_22_0": value  <=  1;
            "HEIGHT_9_22_1": value  <=  1;
            "HEIGHT_9_23_0": value  <=  6;
            "HEIGHT_9_23_1": value  <=  2;
            "HEIGHT_9_24_0": value  <=  2;
            "HEIGHT_9_24_1": value  <=  2;
            "HEIGHT_9_25_0": value  <=  3;
            "HEIGHT_9_25_1": value  <=  1;
            "HEIGHT_9_26_0": value  <=  3;
            "HEIGHT_9_26_1": value  <=  1;
            "HEIGHT_9_27_0": value  <=  2;
            "HEIGHT_9_27_1": value  <=  1;
            "HEIGHT_9_28_0": value  <=  3;
            "HEIGHT_9_28_1": value  <=  1;
            "HEIGHT_9_29_0": value  <=  6;
            "HEIGHT_9_29_1": value  <=  2;
            "HEIGHT_9_30_0": value  <=  6;
            "HEIGHT_9_30_1": value  <=  2;
            "HEIGHT_9_31_0": value  <=  9;
            "HEIGHT_9_31_1": value  <=  3;
            "HEIGHT_9_32_0": value  <=  6;
            "HEIGHT_9_32_1": value  <=  2;
            "HEIGHT_9_33_0": value  <=  2;
            "HEIGHT_9_33_1": value  <=  2;
            "HEIGHT_9_34_0": value  <=  2;
            "HEIGHT_9_34_1": value  <=  2;
            "HEIGHT_9_35_0": value  <=  6;
            "HEIGHT_9_35_1": value  <=  2;
            "HEIGHT_9_36_0": value  <=  6;
            "HEIGHT_9_36_1": value  <=  2;
            "HEIGHT_9_37_0": value  <=  3;
            "HEIGHT_9_37_1": value  <=  1;
            "HEIGHT_9_38_0": value  <=  9;
            "HEIGHT_9_38_1": value  <=  3;
            "HEIGHT_9_39_0": value  <=  15;
            "HEIGHT_9_39_1": value  <=  15;
            "HEIGHT_9_40_0": value  <=  2;
            "HEIGHT_9_40_1": value  <=  1;
            "HEIGHT_9_41_0": value  <=  10;
            "HEIGHT_9_41_1": value  <=  5;
            "HEIGHT_9_42_0": value  <=  12;
            "HEIGHT_9_42_1": value  <=  12;
            "HEIGHT_9_43_0": value  <=  2;
            "HEIGHT_9_43_1": value  <=  2;
            "HEIGHT_9_44_0": value  <=  2;
            "HEIGHT_9_44_1": value  <=  2;
            "HEIGHT_9_45_0": value  <=  5;
            "HEIGHT_9_45_1": value  <=  5;
            "HEIGHT_9_46_0": value  <=  10;
            "HEIGHT_9_46_1": value  <=  10;
            "HEIGHT_9_47_0": value  <=  2;
            "HEIGHT_9_47_1": value  <=  2;
            "HEIGHT_9_48_0": value  <=  8;
            "HEIGHT_9_48_1": value  <=  4;
            "HEIGHT_9_49_0": value  <=  3;
            "HEIGHT_9_49_1": value  <=  1;
            "HEIGHT_9_50_0": value  <=  3;
            "HEIGHT_9_50_1": value  <=  1;
            "HEIGHT_9_51_0": value  <=  2;
            "HEIGHT_9_51_1": value  <=  2;
            "HEIGHT_9_52_0": value  <=  4;
            "HEIGHT_9_52_1": value  <=  2;
            "HEIGHT_9_52_2": value  <=  2;
            "HEIGHT_9_53_0": value  <=  4;
            "HEIGHT_9_53_1": value  <=  2;
            "HEIGHT_9_53_2": value  <=  2;
            "HEIGHT_9_54_0": value  <=  12;
            "HEIGHT_9_54_1": value  <=  12;
            "HEIGHT_9_55_0": value  <=  2;
            "HEIGHT_9_55_1": value  <=  2;
            "HEIGHT_9_56_0": value  <=  5;
            "HEIGHT_9_56_1": value  <=  5;
            "HEIGHT_9_57_0": value  <=  4;
            "HEIGHT_9_57_1": value  <=  2;
            "HEIGHT_9_57_2": value  <=  2;
            "HEIGHT_9_58_0": value  <=  2;
            "HEIGHT_9_58_1": value  <=  1;
            "HEIGHT_9_59_0": value  <=  4;
            "HEIGHT_9_59_1": value  <=  2;
            "HEIGHT_9_59_2": value  <=  2;
            "HEIGHT_9_60_0": value  <=  4;
            "HEIGHT_9_60_1": value  <=  2;
            "HEIGHT_9_60_2": value  <=  2;
            "HEIGHT_9_61_0": value  <=  12;
            "HEIGHT_9_61_1": value  <=  6;
            "HEIGHT_9_62_0": value  <=  6;
            "HEIGHT_9_62_1": value  <=  6;
            "HEIGHT_9_63_0": value  <=  3;
            "HEIGHT_9_63_1": value  <=  1;
            "HEIGHT_9_64_0": value  <=  3;
            "HEIGHT_9_64_1": value  <=  1;
            "HEIGHT_9_65_0": value  <=  3;
            "HEIGHT_9_65_1": value  <=  1;
            "HEIGHT_9_66_0": value  <=  4;
            "HEIGHT_9_66_1": value  <=  2;
            "HEIGHT_9_66_2": value  <=  2;
            "HEIGHT_9_67_0": value  <=  3;
            "HEIGHT_9_67_1": value  <=  1;
            "HEIGHT_9_68_0": value  <=  12;
            "HEIGHT_9_68_1": value  <=  6;
            "HEIGHT_9_69_0": value  <=  5;
            "HEIGHT_9_69_1": value  <=  5;
            "HEIGHT_9_70_0": value  <=  12;
            "HEIGHT_9_70_1": value  <=  6;
            "HEIGHT_10_0_0": value  <=  3;
            "HEIGHT_10_0_1": value  <=  3;
            "HEIGHT_10_1_0": value  <=  10;
            "HEIGHT_10_1_1": value  <=  5;
            "HEIGHT_10_1_2": value  <=  5;
            "HEIGHT_10_2_0": value  <=  12;
            "HEIGHT_10_2_1": value  <=  6;
            "HEIGHT_10_2_2": value  <=  6;
            "HEIGHT_10_3_0": value  <=  6;
            "HEIGHT_10_3_1": value  <=  2;
            "HEIGHT_10_4_0": value  <=  2;
            "HEIGHT_10_4_1": value  <=  1;
            "HEIGHT_10_5_0": value  <=  2;
            "HEIGHT_10_5_1": value  <=  2;
            "HEIGHT_10_6_0": value  <=  16;
            "HEIGHT_10_6_1": value  <=  8;
            "HEIGHT_10_7_0": value  <=  8;
            "HEIGHT_10_7_1": value  <=  4;
            "HEIGHT_10_8_0": value  <=  1;
            "HEIGHT_10_8_1": value  <=  1;
            "HEIGHT_10_9_0": value  <=  4;
            "HEIGHT_10_9_1": value  <=  2;
            "HEIGHT_10_10_0": value  <=  8;
            "HEIGHT_10_10_1": value  <=  4;
            "HEIGHT_10_11_0": value  <=  12;
            "HEIGHT_10_11_1": value  <=  6;
            "HEIGHT_10_12_0": value  <=  2;
            "HEIGHT_10_12_1": value  <=  2;
            "HEIGHT_10_13_0": value  <=  6;
            "HEIGHT_10_13_1": value  <=  2;
            "HEIGHT_10_14_0": value  <=  2;
            "HEIGHT_10_14_1": value  <=  1;
            "HEIGHT_10_15_0": value  <=  3;
            "HEIGHT_10_15_1": value  <=  1;
            "HEIGHT_10_16_0": value  <=  2;
            "HEIGHT_10_16_1": value  <=  1;
            "HEIGHT_10_17_0": value  <=  6;
            "HEIGHT_10_17_1": value  <=  3;
            "HEIGHT_10_17_2": value  <=  3;
            "HEIGHT_10_18_0": value  <=  4;
            "HEIGHT_10_18_1": value  <=  4;
            "HEIGHT_10_19_0": value  <=  3;
            "HEIGHT_10_19_1": value  <=  1;
            "HEIGHT_10_20_0": value  <=  6;
            "HEIGHT_10_20_1": value  <=  2;
            "HEIGHT_10_21_0": value  <=  3;
            "HEIGHT_10_21_1": value  <=  3;
            "HEIGHT_10_22_0": value  <=  14;
            "HEIGHT_10_22_1": value  <=  14;
            "HEIGHT_10_23_0": value  <=  3;
            "HEIGHT_10_23_1": value  <=  3;
            "HEIGHT_10_24_0": value  <=  4;
            "HEIGHT_10_24_1": value  <=  2;
            "HEIGHT_10_25_0": value  <=  6;
            "HEIGHT_10_25_1": value  <=  2;
            "HEIGHT_10_26_0": value  <=  2;
            "HEIGHT_10_26_1": value  <=  1;
            "HEIGHT_10_27_0": value  <=  6;
            "HEIGHT_10_27_1": value  <=  6;
            "HEIGHT_10_28_0": value  <=  1;
            "HEIGHT_10_28_1": value  <=  1;
            "HEIGHT_10_29_0": value  <=  6;
            "HEIGHT_10_29_1": value  <=  6;
            "HEIGHT_10_30_0": value  <=  10;
            "HEIGHT_10_30_1": value  <=  5;
            "HEIGHT_10_31_0": value  <=  6;
            "HEIGHT_10_31_1": value  <=  6;
            "HEIGHT_10_32_0": value  <=  6;
            "HEIGHT_10_32_1": value  <=  6;
            "HEIGHT_10_33_0": value  <=  2;
            "HEIGHT_10_33_1": value  <=  1;
            "HEIGHT_10_34_0": value  <=  8;
            "HEIGHT_10_34_1": value  <=  8;
            "HEIGHT_10_35_0": value  <=  4;
            "HEIGHT_10_35_1": value  <=  2;
            "HEIGHT_10_35_2": value  <=  2;
            "HEIGHT_10_36_0": value  <=  2;
            "HEIGHT_10_36_1": value  <=  1;
            "HEIGHT_10_37_0": value  <=  6;
            "HEIGHT_10_37_1": value  <=  3;
            "HEIGHT_10_37_2": value  <=  3;
            "HEIGHT_10_38_0": value  <=  4;
            "HEIGHT_10_38_1": value  <=  4;
            "HEIGHT_10_39_0": value  <=  3;
            "HEIGHT_10_39_1": value  <=  3;
            "HEIGHT_10_40_0": value  <=  8;
            "HEIGHT_10_40_1": value  <=  8;
            "HEIGHT_10_41_0": value  <=  3;
            "HEIGHT_10_41_1": value  <=  1;
            "HEIGHT_10_42_0": value  <=  1;
            "HEIGHT_10_42_1": value  <=  1;
            "HEIGHT_10_43_0": value  <=  3;
            "HEIGHT_10_43_1": value  <=  1;
            "HEIGHT_10_44_0": value  <=  3;
            "HEIGHT_10_44_1": value  <=  1;
            "HEIGHT_10_45_0": value  <=  2;
            "HEIGHT_10_45_1": value  <=  1;
            "HEIGHT_10_46_0": value  <=  4;
            "HEIGHT_10_46_1": value  <=  2;
            "HEIGHT_10_47_0": value  <=  4;
            "HEIGHT_10_47_1": value  <=  4;
            "HEIGHT_10_48_0": value  <=  3;
            "HEIGHT_10_48_1": value  <=  1;
            "HEIGHT_10_49_0": value  <=  6;
            "HEIGHT_10_49_1": value  <=  2;
            "HEIGHT_10_50_0": value  <=  6;
            "HEIGHT_10_50_1": value  <=  3;
            "HEIGHT_10_51_0": value  <=  6;
            "HEIGHT_10_51_1": value  <=  3;
            "HEIGHT_10_52_0": value  <=  4;
            "HEIGHT_10_52_1": value  <=  4;
            "HEIGHT_10_53_0": value  <=  2;
            "HEIGHT_10_53_1": value  <=  2;
            "HEIGHT_10_54_0": value  <=  4;
            "HEIGHT_10_54_1": value  <=  4;
            "HEIGHT_10_55_0": value  <=  3;
            "HEIGHT_10_55_1": value  <=  3;
            "HEIGHT_10_56_0": value  <=  3;
            "HEIGHT_10_56_1": value  <=  1;
            "HEIGHT_10_57_0": value  <=  12;
            "HEIGHT_10_57_1": value  <=  4;
            "HEIGHT_10_58_0": value  <=  6;
            "HEIGHT_10_58_1": value  <=  3;
            "HEIGHT_10_58_2": value  <=  3;
            "HEIGHT_10_59_0": value  <=  2;
            "HEIGHT_10_59_1": value  <=  1;
            "HEIGHT_10_60_0": value  <=  2;
            "HEIGHT_10_60_1": value  <=  1;
            "HEIGHT_10_61_0": value  <=  3;
            "HEIGHT_10_61_1": value  <=  1;
            "HEIGHT_10_62_0": value  <=  1;
            "HEIGHT_10_62_1": value  <=  1;
            "HEIGHT_10_63_0": value  <=  3;
            "HEIGHT_10_63_1": value  <=  3;
            "HEIGHT_10_64_0": value  <=  2;
            "HEIGHT_10_64_1": value  <=  2;
            "HEIGHT_10_65_0": value  <=  5;
            "HEIGHT_10_65_1": value  <=  5;
            "HEIGHT_10_66_0": value  <=  5;
            "HEIGHT_10_66_1": value  <=  5;
            "HEIGHT_10_67_0": value  <=  5;
            "HEIGHT_10_67_1": value  <=  5;
            "HEIGHT_10_68_0": value  <=  6;
            "HEIGHT_10_68_1": value  <=  6;
            "HEIGHT_10_69_0": value  <=  5;
            "HEIGHT_10_69_1": value  <=  5;
            "HEIGHT_10_70_0": value  <=  2;
            "HEIGHT_10_70_1": value  <=  1;
            "HEIGHT_10_71_0": value  <=  3;
            "HEIGHT_10_71_1": value  <=  1;
            "HEIGHT_10_72_0": value  <=  2;
            "HEIGHT_10_72_1": value  <=  1;
            "HEIGHT_10_72_2": value  <=  1;
            "HEIGHT_10_73_0": value  <=  4;
            "HEIGHT_10_73_1": value  <=  2;
            "HEIGHT_10_73_2": value  <=  2;
            "HEIGHT_10_74_0": value  <=  2;
            "HEIGHT_10_74_1": value  <=  1;
            "HEIGHT_10_74_2": value  <=  1;
            "HEIGHT_10_75_0": value  <=  2;
            "HEIGHT_10_75_1": value  <=  1;
            "HEIGHT_10_76_0": value  <=  3;
            "HEIGHT_10_76_1": value  <=  1;
            "HEIGHT_10_77_0": value  <=  3;
            "HEIGHT_10_77_1": value  <=  1;
            "HEIGHT_10_78_0": value  <=  3;
            "HEIGHT_10_78_1": value  <=  1;
            "HEIGHT_10_79_0": value  <=  3;
            "HEIGHT_10_79_1": value  <=  1;
            "HEIGHT_11_0_0": value  <=  4;
            "HEIGHT_11_0_1": value  <=  2;
            "HEIGHT_11_1_0": value  <=  4;
            "HEIGHT_11_1_1": value  <=  2;
            "HEIGHT_11_1_2": value  <=  2;
            "HEIGHT_11_2_0": value  <=  6;
            "HEIGHT_11_2_1": value  <=  2;
            "HEIGHT_11_3_0": value  <=  4;
            "HEIGHT_11_3_1": value  <=  2;
            "HEIGHT_11_3_2": value  <=  2;
            "HEIGHT_11_4_0": value  <=  2;
            "HEIGHT_11_4_1": value  <=  1;
            "HEIGHT_11_5_0": value  <=  3;
            "HEIGHT_11_5_1": value  <=  3;
            "HEIGHT_11_6_0": value  <=  4;
            "HEIGHT_11_6_1": value  <=  2;
            "HEIGHT_11_6_2": value  <=  2;
            "HEIGHT_11_7_0": value  <=  7;
            "HEIGHT_11_7_1": value  <=  7;
            "HEIGHT_11_8_0": value  <=  3;
            "HEIGHT_11_8_1": value  <=  3;
            "HEIGHT_11_9_0": value  <=  2;
            "HEIGHT_11_9_1": value  <=  1;
            "HEIGHT_11_10_0": value  <=  3;
            "HEIGHT_11_10_1": value  <=  1;
            "HEIGHT_11_11_0": value  <=  3;
            "HEIGHT_11_11_1": value  <=  3;
            "HEIGHT_11_12_0": value  <=  10;
            "HEIGHT_11_12_1": value  <=  5;
            "HEIGHT_11_13_0": value  <=  2;
            "HEIGHT_11_13_1": value  <=  2;
            "HEIGHT_11_14_0": value  <=  2;
            "HEIGHT_11_14_1": value  <=  2;
            "HEIGHT_11_15_0": value  <=  1;
            "HEIGHT_11_15_1": value  <=  1;
            "HEIGHT_11_16_0": value  <=  2;
            "HEIGHT_11_16_1": value  <=  2;
            "HEIGHT_11_17_0": value  <=  5;
            "HEIGHT_11_17_1": value  <=  5;
            "HEIGHT_11_18_0": value  <=  12;
            "HEIGHT_11_18_1": value  <=  6;
            "HEIGHT_11_19_0": value  <=  3;
            "HEIGHT_11_19_1": value  <=  1;
            "HEIGHT_11_20_0": value  <=  3;
            "HEIGHT_11_20_1": value  <=  3;
            "HEIGHT_11_21_0": value  <=  6;
            "HEIGHT_11_21_1": value  <=  2;
            "HEIGHT_11_22_0": value  <=  6;
            "HEIGHT_11_22_1": value  <=  2;
            "HEIGHT_11_23_0": value  <=  3;
            "HEIGHT_11_23_1": value  <=  1;
            "HEIGHT_11_24_0": value  <=  3;
            "HEIGHT_11_24_1": value  <=  1;
            "HEIGHT_11_25_0": value  <=  6;
            "HEIGHT_11_25_1": value  <=  2;
            "HEIGHT_11_26_0": value  <=  6;
            "HEIGHT_11_26_1": value  <=  2;
            "HEIGHT_11_27_0": value  <=  3;
            "HEIGHT_11_27_1": value  <=  1;
            "HEIGHT_11_28_0": value  <=  4;
            "HEIGHT_11_28_1": value  <=  4;
            "HEIGHT_11_29_0": value  <=  6;
            "HEIGHT_11_29_1": value  <=  2;
            "HEIGHT_11_30_0": value  <=  2;
            "HEIGHT_11_30_1": value  <=  2;
            "HEIGHT_11_31_0": value  <=  4;
            "HEIGHT_11_31_1": value  <=  2;
            "HEIGHT_11_31_2": value  <=  2;
            "HEIGHT_11_32_0": value  <=  2;
            "HEIGHT_11_32_1": value  <=  1;
            "HEIGHT_11_32_2": value  <=  1;
            "HEIGHT_11_33_0": value  <=  2;
            "HEIGHT_11_33_1": value  <=  1;
            "HEIGHT_11_34_0": value  <=  8;
            "HEIGHT_11_34_1": value  <=  4;
            "HEIGHT_11_35_0": value  <=  2;
            "HEIGHT_11_35_1": value  <=  1;
            "HEIGHT_11_36_0": value  <=  2;
            "HEIGHT_11_36_1": value  <=  1;
            "HEIGHT_11_37_0": value  <=  5;
            "HEIGHT_11_37_1": value  <=  5;
            "HEIGHT_11_38_0": value  <=  8;
            "HEIGHT_11_38_1": value  <=  8;
            "HEIGHT_11_39_0": value  <=  4;
            "HEIGHT_11_39_1": value  <=  4;
            "HEIGHT_11_40_0": value  <=  2;
            "HEIGHT_11_40_1": value  <=  1;
            "HEIGHT_11_41_0": value  <=  3;
            "HEIGHT_11_41_1": value  <=  3;
            "HEIGHT_11_42_0": value  <=  3;
            "HEIGHT_11_42_1": value  <=  3;
            "HEIGHT_11_43_0": value  <=  2;
            "HEIGHT_11_43_1": value  <=  1;
            "HEIGHT_11_44_0": value  <=  9;
            "HEIGHT_11_44_1": value  <=  9;
            "HEIGHT_11_45_0": value  <=  13;
            "HEIGHT_11_45_1": value  <=  13;
            "HEIGHT_11_46_0": value  <=  8;
            "HEIGHT_11_46_1": value  <=  4;
            "HEIGHT_11_46_2": value  <=  4;
            "HEIGHT_11_47_0": value  <=  11;
            "HEIGHT_11_47_1": value  <=  11;
            "HEIGHT_11_48_0": value  <=  12;
            "HEIGHT_11_48_1": value  <=  6;
            "HEIGHT_11_48_2": value  <=  6;
            "HEIGHT_11_49_0": value  <=  3;
            "HEIGHT_11_49_1": value  <=  1;
            "HEIGHT_11_50_0": value  <=  2;
            "HEIGHT_11_50_1": value  <=  1;
            "HEIGHT_11_51_0": value  <=  2;
            "HEIGHT_11_51_1": value  <=  2;
            "HEIGHT_11_52_0": value  <=  2;
            "HEIGHT_11_52_1": value  <=  2;
            "HEIGHT_11_53_0": value  <=  2;
            "HEIGHT_11_53_1": value  <=  2;
            "HEIGHT_11_54_0": value  <=  3;
            "HEIGHT_11_54_1": value  <=  1;
            "HEIGHT_11_55_0": value  <=  3;
            "HEIGHT_11_55_1": value  <=  3;
            "HEIGHT_11_56_0": value  <=  2;
            "HEIGHT_11_56_1": value  <=  1;
            "HEIGHT_11_56_2": value  <=  1;
            "HEIGHT_11_57_0": value  <=  3;
            "HEIGHT_11_57_1": value  <=  1;
            "HEIGHT_11_58_0": value  <=  2;
            "HEIGHT_11_58_1": value  <=  1;
            "HEIGHT_11_59_0": value  <=  2;
            "HEIGHT_11_59_1": value  <=  1;
            "HEIGHT_11_60_0": value  <=  4;
            "HEIGHT_11_60_1": value  <=  2;
            "HEIGHT_11_60_2": value  <=  2;
            "HEIGHT_11_61_0": value  <=  3;
            "HEIGHT_11_61_1": value  <=  1;
            "HEIGHT_11_62_0": value  <=  3;
            "HEIGHT_11_62_1": value  <=  1;
            "HEIGHT_11_63_0": value  <=  3;
            "HEIGHT_11_63_1": value  <=  1;
            "HEIGHT_11_64_0": value  <=  3;
            "HEIGHT_11_64_1": value  <=  1;
            "HEIGHT_11_65_0": value  <=  2;
            "HEIGHT_11_65_1": value  <=  1;
            "HEIGHT_11_66_0": value  <=  2;
            "HEIGHT_11_66_1": value  <=  1;
            "HEIGHT_11_67_0": value  <=  3;
            "HEIGHT_11_67_1": value  <=  1;
            "HEIGHT_11_68_0": value  <=  3;
            "HEIGHT_11_68_1": value  <=  3;
            "HEIGHT_11_69_0": value  <=  2;
            "HEIGHT_11_69_1": value  <=  1;
            "HEIGHT_11_70_0": value  <=  2;
            "HEIGHT_11_70_1": value  <=  2;
            "HEIGHT_11_71_0": value  <=  2;
            "HEIGHT_11_71_1": value  <=  1;
            "HEIGHT_11_72_0": value  <=  2;
            "HEIGHT_11_72_1": value  <=  1;
            "HEIGHT_11_73_0": value  <=  3;
            "HEIGHT_11_73_1": value  <=  1;
            "HEIGHT_11_74_0": value  <=  3;
            "HEIGHT_11_74_1": value  <=  1;
            "HEIGHT_11_75_0": value  <=  14;
            "HEIGHT_11_75_1": value  <=  14;
            "HEIGHT_11_76_0": value  <=  14;
            "HEIGHT_11_76_1": value  <=  14;
            "HEIGHT_11_77_0": value  <=  3;
            "HEIGHT_11_77_1": value  <=  1;
            "HEIGHT_11_78_0": value  <=  1;
            "HEIGHT_11_78_1": value  <=  1;
            "HEIGHT_11_79_0": value  <=  3;
            "HEIGHT_11_79_1": value  <=  1;
            "HEIGHT_11_80_0": value  <=  3;
            "HEIGHT_11_80_1": value  <=  3;
            "HEIGHT_11_81_0": value  <=  18;
            "HEIGHT_11_81_1": value  <=  9;
            "HEIGHT_11_82_0": value  <=  14;
            "HEIGHT_11_82_1": value  <=  7;
            "HEIGHT_11_83_0": value  <=  4;
            "HEIGHT_11_83_1": value  <=  4;
            "HEIGHT_11_84_0": value  <=  3;
            "HEIGHT_11_84_1": value  <=  1;
            "HEIGHT_11_85_0": value  <=  3;
            "HEIGHT_11_85_1": value  <=  1;
            "HEIGHT_11_86_0": value  <=  14;
            "HEIGHT_11_86_1": value  <=  7;
            "HEIGHT_11_86_2": value  <=  7;
            "HEIGHT_11_87_0": value  <=  18;
            "HEIGHT_11_87_1": value  <=  9;
            "HEIGHT_11_87_2": value  <=  9;
            "HEIGHT_11_88_0": value  <=  3;
            "HEIGHT_11_88_1": value  <=  1;
            "HEIGHT_11_89_0": value  <=  18;
            "HEIGHT_11_89_1": value  <=  9;
            "HEIGHT_11_89_2": value  <=  9;
            "HEIGHT_11_90_0": value  <=  3;
            "HEIGHT_11_90_1": value  <=  1;
            "HEIGHT_11_91_0": value  <=  3;
            "HEIGHT_11_91_1": value  <=  1;
            "HEIGHT_11_92_0": value  <=  9;
            "HEIGHT_11_92_1": value  <=  3;
            "HEIGHT_11_93_0": value  <=  11;
            "HEIGHT_11_93_1": value  <=  11;
            "HEIGHT_11_94_0": value  <=  1;
            "HEIGHT_11_94_1": value  <=  1;
            "HEIGHT_11_95_0": value  <=  7;
            "HEIGHT_11_95_1": value  <=  7;
            "HEIGHT_11_96_0": value  <=  7;
            "HEIGHT_11_96_1": value  <=  7;
            "HEIGHT_11_97_0": value  <=  12;
            "HEIGHT_11_97_1": value  <=  4;
            "HEIGHT_11_98_0": value  <=  11;
            "HEIGHT_11_98_1": value  <=  11;
            "HEIGHT_11_99_0": value  <=  20;
            "HEIGHT_11_99_1": value  <=  20;
            "HEIGHT_11_100_0": value  <=  2;
            "HEIGHT_11_100_1": value  <=  1;
            "HEIGHT_11_101_0": value  <=  8;
            "HEIGHT_11_101_1": value  <=  4;
            "HEIGHT_11_101_2": value  <=  4;
            "HEIGHT_11_102_0": value  <=  4;
            "HEIGHT_11_102_1": value  <=  2;
            "HEIGHT_11_102_2": value  <=  2;
            "HEIGHT_12_0_0": value  <=  4;
            "HEIGHT_12_0_1": value  <=  4;
            "HEIGHT_12_1_0": value  <=  4;
            "HEIGHT_12_1_1": value  <=  2;
            "HEIGHT_12_1_2": value  <=  2;
            "HEIGHT_12_2_0": value  <=  6;
            "HEIGHT_12_2_1": value  <=  3;
            "HEIGHT_12_3_0": value  <=  4;
            "HEIGHT_12_3_1": value  <=  2;
            "HEIGHT_12_3_2": value  <=  2;
            "HEIGHT_12_4_0": value  <=  12;
            "HEIGHT_12_4_1": value  <=  6;
            "HEIGHT_12_5_0": value  <=  18;
            "HEIGHT_12_5_1": value  <=  18;
            "HEIGHT_12_6_0": value  <=  2;
            "HEIGHT_12_6_1": value  <=  2;
            "HEIGHT_12_7_0": value  <=  2;
            "HEIGHT_12_7_1": value  <=  1;
            "HEIGHT_12_8_0": value  <=  6;
            "HEIGHT_12_8_1": value  <=  6;
            "HEIGHT_12_9_0": value  <=  2;
            "HEIGHT_12_9_1": value  <=  1;
            "HEIGHT_12_10_0": value  <=  4;
            "HEIGHT_12_10_1": value  <=  2;
            "HEIGHT_12_11_0": value  <=  12;
            "HEIGHT_12_11_1": value  <=  12;
            "HEIGHT_12_12_0": value  <=  3;
            "HEIGHT_12_12_1": value  <=  1;
            "HEIGHT_12_13_0": value  <=  17;
            "HEIGHT_12_13_1": value  <=  17;
            "HEIGHT_12_14_0": value  <=  1;
            "HEIGHT_12_14_1": value  <=  1;
            "HEIGHT_12_15_0": value  <=  3;
            "HEIGHT_12_15_1": value  <=  1;
            "HEIGHT_12_16_0": value  <=  4;
            "HEIGHT_12_16_1": value  <=  2;
            "HEIGHT_12_17_0": value  <=  10;
            "HEIGHT_12_17_1": value  <=  5;
            "HEIGHT_12_18_0": value  <=  2;
            "HEIGHT_12_18_1": value  <=  2;
            "HEIGHT_12_19_0": value  <=  6;
            "HEIGHT_12_19_1": value  <=  2;
            "HEIGHT_12_20_0": value  <=  6;
            "HEIGHT_12_20_1": value  <=  6;
            "HEIGHT_12_21_0": value  <=  6;
            "HEIGHT_12_21_1": value  <=  2;
            "HEIGHT_12_22_0": value  <=  4;
            "HEIGHT_12_22_1": value  <=  4;
            "HEIGHT_12_23_0": value  <=  3;
            "HEIGHT_12_23_1": value  <=  1;
            "HEIGHT_12_24_0": value  <=  3;
            "HEIGHT_12_24_1": value  <=  1;
            "HEIGHT_12_25_0": value  <=  3;
            "HEIGHT_12_25_1": value  <=  1;
            "HEIGHT_12_26_0": value  <=  3;
            "HEIGHT_12_26_1": value  <=  1;
            "HEIGHT_12_27_0": value  <=  7;
            "HEIGHT_12_27_1": value  <=  7;
            "HEIGHT_12_28_0": value  <=  6;
            "HEIGHT_12_28_1": value  <=  2;
            "HEIGHT_12_29_0": value  <=  3;
            "HEIGHT_12_29_1": value  <=  1;
            "HEIGHT_12_30_0": value  <=  14;
            "HEIGHT_12_30_1": value  <=  14;
            "HEIGHT_12_31_0": value  <=  6;
            "HEIGHT_12_31_1": value  <=  2;
            "HEIGHT_12_32_0": value  <=  6;
            "HEIGHT_12_32_1": value  <=  2;
            "HEIGHT_12_33_0": value  <=  2;
            "HEIGHT_12_33_1": value  <=  1;
            "HEIGHT_12_33_2": value  <=  1;
            "HEIGHT_12_34_0": value  <=  14;
            "HEIGHT_12_34_1": value  <=  14;
            "HEIGHT_12_35_0": value  <=  3;
            "HEIGHT_12_35_1": value  <=  1;
            "HEIGHT_12_36_0": value  <=  3;
            "HEIGHT_12_36_1": value  <=  1;
            "HEIGHT_12_37_0": value  <=  6;
            "HEIGHT_12_37_1": value  <=  3;
            "HEIGHT_12_38_0": value  <=  9;
            "HEIGHT_12_38_1": value  <=  3;
            "HEIGHT_12_39_0": value  <=  2;
            "HEIGHT_12_39_1": value  <=  1;
            "HEIGHT_12_39_2": value  <=  1;
            "HEIGHT_12_40_0": value  <=  3;
            "HEIGHT_12_40_1": value  <=  1;
            "HEIGHT_12_41_0": value  <=  3;
            "HEIGHT_12_41_1": value  <=  1;
            "HEIGHT_12_42_0": value  <=  6;
            "HEIGHT_12_42_1": value  <=  6;
            "HEIGHT_12_43_0": value  <=  6;
            "HEIGHT_12_43_1": value  <=  6;
            "HEIGHT_12_44_0": value  <=  3;
            "HEIGHT_12_44_1": value  <=  1;
            "HEIGHT_12_45_0": value  <=  3;
            "HEIGHT_12_45_1": value  <=  1;
            "HEIGHT_12_46_0": value  <=  3;
            "HEIGHT_12_46_1": value  <=  1;
            "HEIGHT_12_47_0": value  <=  12;
            "HEIGHT_12_47_1": value  <=  6;
            "HEIGHT_12_48_0": value  <=  10;
            "HEIGHT_12_48_1": value  <=  5;
            "HEIGHT_12_48_2": value  <=  5;
            "HEIGHT_12_49_0": value  <=  3;
            "HEIGHT_12_49_1": value  <=  1;
            "HEIGHT_12_50_0": value  <=  3;
            "HEIGHT_12_50_1": value  <=  1;
            "HEIGHT_12_51_0": value  <=  5;
            "HEIGHT_12_51_1": value  <=  5;
            "HEIGHT_12_52_0": value  <=  6;
            "HEIGHT_12_52_1": value  <=  2;
            "HEIGHT_12_53_0": value  <=  2;
            "HEIGHT_12_53_1": value  <=  1;
            "HEIGHT_12_54_0": value  <=  1;
            "HEIGHT_12_54_1": value  <=  1;
            "HEIGHT_12_55_0": value  <=  2;
            "HEIGHT_12_55_1": value  <=  1;
            "HEIGHT_12_55_2": value  <=  1;
            "HEIGHT_12_56_0": value  <=  2;
            "HEIGHT_12_56_1": value  <=  1;
            "HEIGHT_12_56_2": value  <=  1;
            "HEIGHT_12_57_0": value  <=  4;
            "HEIGHT_12_57_1": value  <=  2;
            "HEIGHT_12_58_0": value  <=  8;
            "HEIGHT_12_58_1": value  <=  8;
            "HEIGHT_12_59_0": value  <=  3;
            "HEIGHT_12_59_1": value  <=  1;
            "HEIGHT_12_60_0": value  <=  4;
            "HEIGHT_12_60_1": value  <=  4;
            "HEIGHT_12_61_0": value  <=  10;
            "HEIGHT_12_61_1": value  <=  5;
            "HEIGHT_12_61_2": value  <=  5;
            "HEIGHT_12_62_0": value  <=  2;
            "HEIGHT_12_62_1": value  <=  1;
            "HEIGHT_12_62_2": value  <=  1;
            "HEIGHT_12_63_0": value  <=  8;
            "HEIGHT_12_63_1": value  <=  8;
            "HEIGHT_12_64_0": value  <=  8;
            "HEIGHT_12_64_1": value  <=  8;
            "HEIGHT_12_65_0": value  <=  7;
            "HEIGHT_12_65_1": value  <=  7;
            "HEIGHT_12_66_0": value  <=  1;
            "HEIGHT_12_66_1": value  <=  1;
            "HEIGHT_12_67_0": value  <=  3;
            "HEIGHT_12_67_1": value  <=  1;
            "HEIGHT_12_68_0": value  <=  2;
            "HEIGHT_12_68_1": value  <=  1;
            "HEIGHT_12_68_2": value  <=  1;
            "HEIGHT_12_69_0": value  <=  3;
            "HEIGHT_12_69_1": value  <=  1;
            "HEIGHT_12_70_0": value  <=  7;
            "HEIGHT_12_70_1": value  <=  7;
            "HEIGHT_12_71_0": value  <=  7;
            "HEIGHT_12_71_1": value  <=  7;
            "HEIGHT_12_72_0": value  <=  20;
            "HEIGHT_12_72_1": value  <=  10;
            "HEIGHT_12_73_0": value  <=  6;
            "HEIGHT_12_73_1": value  <=  2;
            "HEIGHT_12_74_0": value  <=  2;
            "HEIGHT_12_74_1": value  <=  1;
            "HEIGHT_12_75_0": value  <=  5;
            "HEIGHT_12_75_1": value  <=  5;
            "HEIGHT_12_76_0": value  <=  4;
            "HEIGHT_12_76_1": value  <=  4;
            "HEIGHT_12_77_0": value  <=  5;
            "HEIGHT_12_77_1": value  <=  5;
            "HEIGHT_12_78_0": value  <=  13;
            "HEIGHT_12_78_1": value  <=  13;
            "HEIGHT_12_79_0": value  <=  5;
            "HEIGHT_12_79_1": value  <=  5;
            "HEIGHT_12_80_0": value  <=  5;
            "HEIGHT_12_80_1": value  <=  5;
            "HEIGHT_12_81_0": value  <=  6;
            "HEIGHT_12_81_1": value  <=  2;
            "HEIGHT_12_82_0": value  <=  6;
            "HEIGHT_12_82_1": value  <=  2;
            "HEIGHT_12_83_0": value  <=  3;
            "HEIGHT_12_83_1": value  <=  1;
            "HEIGHT_12_84_0": value  <=  10;
            "HEIGHT_12_84_1": value  <=  5;
            "HEIGHT_12_84_2": value  <=  5;
            "HEIGHT_12_85_0": value  <=  4;
            "HEIGHT_12_85_1": value  <=  2;
            "HEIGHT_12_86_0": value  <=  3;
            "HEIGHT_12_86_1": value  <=  1;
            "HEIGHT_12_87_0": value  <=  3;
            "HEIGHT_12_87_1": value  <=  1;
            "HEIGHT_12_88_0": value  <=  5;
            "HEIGHT_12_88_1": value  <=  5;
            "HEIGHT_12_89_0": value  <=  5;
            "HEIGHT_12_89_1": value  <=  5;
            "HEIGHT_12_90_0": value  <=  5;
            "HEIGHT_12_90_1": value  <=  5;
            "HEIGHT_12_91_0": value  <=  14;
            "HEIGHT_12_91_1": value  <=  14;
            "HEIGHT_12_92_0": value  <=  6;
            "HEIGHT_12_92_1": value  <=  2;
            "HEIGHT_12_93_0": value  <=  4;
            "HEIGHT_12_93_1": value  <=  4;
            "HEIGHT_12_94_0": value  <=  10;
            "HEIGHT_12_94_1": value  <=  10;
            "HEIGHT_12_95_0": value  <=  14;
            "HEIGHT_12_95_1": value  <=  14;
            "HEIGHT_12_96_0": value  <=  14;
            "HEIGHT_12_96_1": value  <=  14;
            "HEIGHT_12_97_0": value  <=  3;
            "HEIGHT_12_97_1": value  <=  1;
            "HEIGHT_12_98_0": value  <=  3;
            "HEIGHT_12_98_1": value  <=  3;
            "HEIGHT_12_99_0": value  <=  18;
            "HEIGHT_12_99_1": value  <=  9;
            "HEIGHT_12_99_2": value  <=  9;
            "HEIGHT_12_100_0": value  <=  3;
            "HEIGHT_12_100_1": value  <=  1;
            "HEIGHT_12_101_0": value  <=  18;
            "HEIGHT_12_101_1": value  <=  9;
            "HEIGHT_12_101_2": value  <=  9;
            "HEIGHT_12_102_0": value  <=  6;
            "HEIGHT_12_102_1": value  <=  3;
            "HEIGHT_12_102_2": value  <=  3;
            "HEIGHT_12_103_0": value  <=  6;
            "HEIGHT_12_103_1": value  <=  2;
            "HEIGHT_12_104_0": value  <=  10;
            "HEIGHT_12_104_1": value  <=  5;
            "HEIGHT_12_104_2": value  <=  5;
            "HEIGHT_12_105_0": value  <=  4;
            "HEIGHT_12_105_1": value  <=  4;
            "HEIGHT_12_106_0": value  <=  6;
            "HEIGHT_12_106_1": value  <=  3;
            "HEIGHT_12_107_0": value  <=  8;
            "HEIGHT_12_107_1": value  <=  4;
            "HEIGHT_12_108_0": value  <=  6;
            "HEIGHT_12_108_1": value  <=  3;
            "HEIGHT_12_108_2": value  <=  3;
            "HEIGHT_12_109_0": value  <=  2;
            "HEIGHT_12_109_1": value  <=  2;
            "HEIGHT_12_110_0": value  <=  5;
            "HEIGHT_12_110_1": value  <=  5;
            "HEIGHT_13_0_0": value  <=  3;
            "HEIGHT_13_0_1": value  <=  3;
            "HEIGHT_13_1_0": value  <=  4;
            "HEIGHT_13_1_1": value  <=  4;
            "HEIGHT_13_2_0": value  <=  4;
            "HEIGHT_13_2_1": value  <=  2;
            "HEIGHT_13_3_0": value  <=  9;
            "HEIGHT_13_3_1": value  <=  3;
            "HEIGHT_13_4_0": value  <=  6;
            "HEIGHT_13_4_1": value  <=  2;
            "HEIGHT_13_5_0": value  <=  4;
            "HEIGHT_13_5_1": value  <=  2;
            "HEIGHT_13_5_2": value  <=  2;
            "HEIGHT_13_6_0": value  <=  4;
            "HEIGHT_13_6_1": value  <=  2;
            "HEIGHT_13_6_2": value  <=  2;
            "HEIGHT_13_7_0": value  <=  8;
            "HEIGHT_13_7_1": value  <=  4;
            "HEIGHT_13_8_0": value  <=  12;
            "HEIGHT_13_8_1": value  <=  6;
            "HEIGHT_13_9_0": value  <=  12;
            "HEIGHT_13_9_1": value  <=  6;
            "HEIGHT_13_9_2": value  <=  6;
            "HEIGHT_13_10_0": value  <=  3;
            "HEIGHT_13_10_1": value  <=  1;
            "HEIGHT_13_11_0": value  <=  5;
            "HEIGHT_13_11_1": value  <=  5;
            "HEIGHT_13_12_0": value  <=  4;
            "HEIGHT_13_12_1": value  <=  2;
            "HEIGHT_13_13_0": value  <=  5;
            "HEIGHT_13_13_1": value  <=  5;
            "HEIGHT_13_14_0": value  <=  5;
            "HEIGHT_13_14_1": value  <=  5;
            "HEIGHT_13_15_0": value  <=  1;
            "HEIGHT_13_15_1": value  <=  1;
            "HEIGHT_13_16_0": value  <=  1;
            "HEIGHT_13_16_1": value  <=  1;
            "HEIGHT_13_17_0": value  <=  3;
            "HEIGHT_13_17_1": value  <=  1;
            "HEIGHT_13_18_0": value  <=  4;
            "HEIGHT_13_18_1": value  <=  2;
            "HEIGHT_13_19_0": value  <=  3;
            "HEIGHT_13_19_1": value  <=  1;
            "HEIGHT_13_20_0": value  <=  2;
            "HEIGHT_13_20_1": value  <=  2;
            "HEIGHT_13_21_0": value  <=  2;
            "HEIGHT_13_21_1": value  <=  1;
            "HEIGHT_13_22_0": value  <=  3;
            "HEIGHT_13_22_1": value  <=  1;
            "HEIGHT_13_23_0": value  <=  4;
            "HEIGHT_13_23_1": value  <=  2;
            "HEIGHT_13_24_0": value  <=  3;
            "HEIGHT_13_24_1": value  <=  1;
            "HEIGHT_13_25_0": value  <=  2;
            "HEIGHT_13_25_1": value  <=  1;
            "HEIGHT_13_26_0": value  <=  9;
            "HEIGHT_13_26_1": value  <=  3;
            "HEIGHT_13_27_0": value  <=  3;
            "HEIGHT_13_27_1": value  <=  1;
            "HEIGHT_13_28_0": value  <=  3;
            "HEIGHT_13_28_1": value  <=  1;
            "HEIGHT_13_29_0": value  <=  6;
            "HEIGHT_13_29_1": value  <=  6;
            "HEIGHT_13_30_0": value  <=  4;
            "HEIGHT_13_30_1": value  <=  4;
            "HEIGHT_13_31_0": value  <=  12;
            "HEIGHT_13_31_1": value  <=  6;
            "HEIGHT_13_31_2": value  <=  6;
            "HEIGHT_13_32_0": value  <=  12;
            "HEIGHT_13_32_1": value  <=  6;
            "HEIGHT_13_32_2": value  <=  6;
            "HEIGHT_13_33_0": value  <=  3;
            "HEIGHT_13_33_1": value  <=  1;
            "HEIGHT_13_34_0": value  <=  2;
            "HEIGHT_13_34_1": value  <=  1;
            "HEIGHT_13_35_0": value  <=  3;
            "HEIGHT_13_35_1": value  <=  1;
            "HEIGHT_13_36_0": value  <=  6;
            "HEIGHT_13_36_1": value  <=  2;
            "HEIGHT_13_37_0": value  <=  3;
            "HEIGHT_13_37_1": value  <=  1;
            "HEIGHT_13_38_0": value  <=  3;
            "HEIGHT_13_38_1": value  <=  1;
            "HEIGHT_13_39_0": value  <=  3;
            "HEIGHT_13_39_1": value  <=  1;
            "HEIGHT_13_40_0": value  <=  3;
            "HEIGHT_13_40_1": value  <=  1;
            "HEIGHT_13_41_0": value  <=  3;
            "HEIGHT_13_41_1": value  <=  1;
            "HEIGHT_13_42_0": value  <=  2;
            "HEIGHT_13_42_1": value  <=  2;
            "HEIGHT_13_43_0": value  <=  3;
            "HEIGHT_13_43_1": value  <=  1;
            "HEIGHT_13_44_0": value  <=  3;
            "HEIGHT_13_44_1": value  <=  1;
            "HEIGHT_13_45_0": value  <=  6;
            "HEIGHT_13_45_1": value  <=  3;
            "HEIGHT_13_45_2": value  <=  3;
            "HEIGHT_13_46_0": value  <=  3;
            "HEIGHT_13_46_1": value  <=  3;
            "HEIGHT_13_47_0": value  <=  4;
            "HEIGHT_13_47_1": value  <=  2;
            "HEIGHT_13_48_0": value  <=  2;
            "HEIGHT_13_48_1": value  <=  1;
            "HEIGHT_13_48_2": value  <=  1;
            "HEIGHT_13_49_0": value  <=  4;
            "HEIGHT_13_49_1": value  <=  4;
            "HEIGHT_13_50_0": value  <=  1;
            "HEIGHT_13_50_1": value  <=  1;
            "HEIGHT_13_51_0": value  <=  2;
            "HEIGHT_13_51_1": value  <=  1;
            "HEIGHT_13_52_0": value  <=  6;
            "HEIGHT_13_52_1": value  <=  2;
            "HEIGHT_13_53_0": value  <=  8;
            "HEIGHT_13_53_1": value  <=  4;
            "HEIGHT_13_53_2": value  <=  4;
            "HEIGHT_13_54_0": value  <=  6;
            "HEIGHT_13_54_1": value  <=  3;
            "HEIGHT_13_54_2": value  <=  3;
            "HEIGHT_13_55_0": value  <=  2;
            "HEIGHT_13_55_1": value  <=  1;
            "HEIGHT_13_56_0": value  <=  3;
            "HEIGHT_13_56_1": value  <=  1;
            "HEIGHT_13_57_0": value  <=  2;
            "HEIGHT_13_57_1": value  <=  1;
            "HEIGHT_13_58_0": value  <=  2;
            "HEIGHT_13_58_1": value  <=  1;
            "HEIGHT_13_59_0": value  <=  2;
            "HEIGHT_13_59_1": value  <=  1;
            "HEIGHT_13_60_0": value  <=  3;
            "HEIGHT_13_60_1": value  <=  1;
            "HEIGHT_13_61_0": value  <=  6;
            "HEIGHT_13_61_1": value  <=  3;
            "HEIGHT_13_62_0": value  <=  12;
            "HEIGHT_13_62_1": value  <=  6;
            "HEIGHT_13_63_0": value  <=  6;
            "HEIGHT_13_63_1": value  <=  3;
            "HEIGHT_13_64_0": value  <=  6;
            "HEIGHT_13_64_1": value  <=  3;
            "HEIGHT_13_65_0": value  <=  3;
            "HEIGHT_13_65_1": value  <=  1;
            "HEIGHT_13_66_0": value  <=  10;
            "HEIGHT_13_66_1": value  <=  5;
            "HEIGHT_13_67_0": value  <=  2;
            "HEIGHT_13_67_1": value  <=  1;
            "HEIGHT_13_68_0": value  <=  3;
            "HEIGHT_13_68_1": value  <=  1;
            "HEIGHT_13_69_0": value  <=  1;
            "HEIGHT_13_69_1": value  <=  1;
            "HEIGHT_13_70_0": value  <=  6;
            "HEIGHT_13_70_1": value  <=  3;
            "HEIGHT_13_70_2": value  <=  3;
            "HEIGHT_13_71_0": value  <=  1;
            "HEIGHT_13_71_1": value  <=  1;
            "HEIGHT_13_72_0": value  <=  1;
            "HEIGHT_13_72_1": value  <=  1;
            "HEIGHT_13_73_0": value  <=  7;
            "HEIGHT_13_73_1": value  <=  7;
            "HEIGHT_13_74_0": value  <=  2;
            "HEIGHT_13_74_1": value  <=  1;
            "HEIGHT_13_75_0": value  <=  9;
            "HEIGHT_13_75_1": value  <=  3;
            "HEIGHT_13_76_0": value  <=  2;
            "HEIGHT_13_76_1": value  <=  2;
            "HEIGHT_13_77_0": value  <=  3;
            "HEIGHT_13_77_1": value  <=  1;
            "HEIGHT_13_78_0": value  <=  3;
            "HEIGHT_13_78_1": value  <=  1;
            "HEIGHT_13_79_0": value  <=  6;
            "HEIGHT_13_79_1": value  <=  6;
            "HEIGHT_13_80_0": value  <=  3;
            "HEIGHT_13_80_1": value  <=  3;
            "HEIGHT_13_81_0": value  <=  6;
            "HEIGHT_13_81_1": value  <=  6;
            "HEIGHT_13_82_0": value  <=  12;
            "HEIGHT_13_82_1": value  <=  6;
            "HEIGHT_13_82_2": value  <=  6;
            "HEIGHT_13_83_0": value  <=  15;
            "HEIGHT_13_83_1": value  <=  15;
            "HEIGHT_13_84_0": value  <=  17;
            "HEIGHT_13_84_1": value  <=  17;
            "HEIGHT_13_85_0": value  <=  7;
            "HEIGHT_13_85_1": value  <=  7;
            "HEIGHT_13_86_0": value  <=  7;
            "HEIGHT_13_86_1": value  <=  7;
            "HEIGHT_13_87_0": value  <=  15;
            "HEIGHT_13_87_1": value  <=  15;
            "HEIGHT_13_88_0": value  <=  15;
            "HEIGHT_13_88_1": value  <=  15;
            "HEIGHT_13_89_0": value  <=  6;
            "HEIGHT_13_89_1": value  <=  2;
            "HEIGHT_13_90_0": value  <=  6;
            "HEIGHT_13_90_1": value  <=  6;
            "HEIGHT_13_91_0": value  <=  6;
            "HEIGHT_13_91_1": value  <=  3;
            "HEIGHT_13_91_2": value  <=  3;
            "HEIGHT_13_92_0": value  <=  9;
            "HEIGHT_13_92_1": value  <=  3;
            "HEIGHT_13_93_0": value  <=  3;
            "HEIGHT_13_93_1": value  <=  1;
            "HEIGHT_13_94_0": value  <=  4;
            "HEIGHT_13_94_1": value  <=  2;
            "HEIGHT_13_95_0": value  <=  12;
            "HEIGHT_13_95_1": value  <=  6;
            "HEIGHT_13_96_0": value  <=  12;
            "HEIGHT_13_96_1": value  <=  6;
            "HEIGHT_13_96_2": value  <=  6;
            "HEIGHT_13_97_0": value  <=  4;
            "HEIGHT_13_97_1": value  <=  2;
            "HEIGHT_13_97_2": value  <=  2;
            "HEIGHT_13_98_0": value  <=  2;
            "HEIGHT_13_98_1": value  <=  1;
            "HEIGHT_13_98_2": value  <=  1;
            "HEIGHT_13_99_0": value  <=  3;
            "HEIGHT_13_99_1": value  <=  1;
            "HEIGHT_13_100_0": value  <=  2;
            "HEIGHT_13_100_1": value  <=  1;
            "HEIGHT_13_101_0": value  <=  2;
            "HEIGHT_13_101_1": value  <=  1;
            "HEIGHT_14_0_0": value  <=  6;
            "HEIGHT_14_0_1": value  <=  2;
            "HEIGHT_14_1_0": value  <=  4;
            "HEIGHT_14_1_1": value  <=  2;
            "HEIGHT_14_1_2": value  <=  2;
            "HEIGHT_14_2_0": value  <=  8;
            "HEIGHT_14_2_1": value  <=  8;
            "HEIGHT_14_3_0": value  <=  12;
            "HEIGHT_14_3_1": value  <=  6;
            "HEIGHT_14_4_0": value  <=  10;
            "HEIGHT_14_4_1": value  <=  5;
            "HEIGHT_14_5_0": value  <=  3;
            "HEIGHT_14_5_1": value  <=  1;
            "HEIGHT_14_6_0": value  <=  6;
            "HEIGHT_14_6_1": value  <=  2;
            "HEIGHT_14_7_0": value  <=  2;
            "HEIGHT_14_7_1": value  <=  1;
            "HEIGHT_14_8_0": value  <=  5;
            "HEIGHT_14_8_1": value  <=  5;
            "HEIGHT_14_9_0": value  <=  6;
            "HEIGHT_14_9_1": value  <=  2;
            "HEIGHT_14_10_0": value  <=  2;
            "HEIGHT_14_10_1": value  <=  1;
            "HEIGHT_14_11_0": value  <=  3;
            "HEIGHT_14_11_1": value  <=  1;
            "HEIGHT_14_12_0": value  <=  6;
            "HEIGHT_14_12_1": value  <=  2;
            "HEIGHT_14_13_0": value  <=  2;
            "HEIGHT_14_13_1": value  <=  1;
            "HEIGHT_14_14_0": value  <=  6;
            "HEIGHT_14_14_1": value  <=  3;
            "HEIGHT_14_14_2": value  <=  3;
            "HEIGHT_14_15_0": value  <=  2;
            "HEIGHT_14_15_1": value  <=  1;
            "HEIGHT_14_16_0": value  <=  12;
            "HEIGHT_14_16_1": value  <=  4;
            "HEIGHT_14_17_0": value  <=  8;
            "HEIGHT_14_17_1": value  <=  4;
            "HEIGHT_14_17_2": value  <=  4;
            "HEIGHT_14_18_0": value  <=  2;
            "HEIGHT_14_18_1": value  <=  2;
            "HEIGHT_14_19_0": value  <=  2;
            "HEIGHT_14_19_1": value  <=  1;
            "HEIGHT_14_20_0": value  <=  12;
            "HEIGHT_14_20_1": value  <=  6;
            "HEIGHT_14_20_2": value  <=  6;
            "HEIGHT_14_21_0": value  <=  10;
            "HEIGHT_14_21_1": value  <=  5;
            "HEIGHT_14_21_2": value  <=  5;
            "HEIGHT_14_22_0": value  <=  6;
            "HEIGHT_14_22_1": value  <=  3;
            "HEIGHT_14_22_2": value  <=  3;
            "HEIGHT_14_23_0": value  <=  10;
            "HEIGHT_14_23_1": value  <=  5;
            "HEIGHT_14_23_2": value  <=  5;
            "HEIGHT_14_24_0": value  <=  2;
            "HEIGHT_14_24_1": value  <=  1;
            "HEIGHT_14_25_0": value  <=  3;
            "HEIGHT_14_25_1": value  <=  1;
            "HEIGHT_14_26_0": value  <=  3;
            "HEIGHT_14_26_1": value  <=  1;
            "HEIGHT_14_27_0": value  <=  4;
            "HEIGHT_14_27_1": value  <=  2;
            "HEIGHT_14_27_2": value  <=  2;
            "HEIGHT_14_28_0": value  <=  3;
            "HEIGHT_14_28_1": value  <=  1;
            "HEIGHT_14_29_0": value  <=  1;
            "HEIGHT_14_29_1": value  <=  1;
            "HEIGHT_14_30_0": value  <=  1;
            "HEIGHT_14_30_1": value  <=  1;
            "HEIGHT_14_31_0": value  <=  15;
            "HEIGHT_14_31_1": value  <=  5;
            "HEIGHT_14_32_0": value  <=  2;
            "HEIGHT_14_32_1": value  <=  2;
            "HEIGHT_14_33_0": value  <=  10;
            "HEIGHT_14_33_1": value  <=  5;
            "HEIGHT_14_33_2": value  <=  5;
            "HEIGHT_14_34_0": value  <=  4;
            "HEIGHT_14_34_1": value  <=  4;
            "HEIGHT_14_35_0": value  <=  8;
            "HEIGHT_14_35_1": value  <=  4;
            "HEIGHT_14_35_2": value  <=  4;
            "HEIGHT_14_36_0": value  <=  3;
            "HEIGHT_14_36_1": value  <=  1;
            "HEIGHT_14_37_0": value  <=  2;
            "HEIGHT_14_37_1": value  <=  2;
            "HEIGHT_14_38_0": value  <=  2;
            "HEIGHT_14_38_1": value  <=  1;
            "HEIGHT_14_39_0": value  <=  14;
            "HEIGHT_14_39_1": value  <=  14;
            "HEIGHT_14_40_0": value  <=  3;
            "HEIGHT_14_40_1": value  <=  3;
            "HEIGHT_14_41_0": value  <=  3;
            "HEIGHT_14_41_1": value  <=  1;
            "HEIGHT_14_42_0": value  <=  6;
            "HEIGHT_14_42_1": value  <=  2;
            "HEIGHT_14_43_0": value  <=  2;
            "HEIGHT_14_43_1": value  <=  1;
            "HEIGHT_14_44_0": value  <=  3;
            "HEIGHT_14_44_1": value  <=  1;
            "HEIGHT_14_45_0": value  <=  9;
            "HEIGHT_14_45_1": value  <=  3;
            "HEIGHT_14_46_0": value  <=  2;
            "HEIGHT_14_46_1": value  <=  2;
            "HEIGHT_14_47_0": value  <=  8;
            "HEIGHT_14_47_1": value  <=  4;
            "HEIGHT_14_47_2": value  <=  4;
            "HEIGHT_14_48_0": value  <=  8;
            "HEIGHT_14_48_1": value  <=  4;
            "HEIGHT_14_48_2": value  <=  4;
            "HEIGHT_14_49_0": value  <=  6;
            "HEIGHT_14_49_1": value  <=  3;
            "HEIGHT_14_49_2": value  <=  3;
            "HEIGHT_14_50_0": value  <=  1;
            "HEIGHT_14_50_1": value  <=  1;
            "HEIGHT_14_51_0": value  <=  6;
            "HEIGHT_14_51_1": value  <=  3;
            "HEIGHT_14_51_2": value  <=  3;
            "HEIGHT_14_52_0": value  <=  3;
            "HEIGHT_14_52_1": value  <=  1;
            "HEIGHT_14_53_0": value  <=  3;
            "HEIGHT_14_53_1": value  <=  1;
            "HEIGHT_14_54_0": value  <=  3;
            "HEIGHT_14_54_1": value  <=  1;
            "HEIGHT_14_55_0": value  <=  6;
            "HEIGHT_14_55_1": value  <=  3;
            "HEIGHT_14_55_2": value  <=  3;
            "HEIGHT_14_56_0": value  <=  6;
            "HEIGHT_14_56_1": value  <=  3;
            "HEIGHT_14_56_2": value  <=  3;
            "HEIGHT_14_57_0": value  <=  2;
            "HEIGHT_14_57_1": value  <=  1;
            "HEIGHT_14_58_0": value  <=  2;
            "HEIGHT_14_58_1": value  <=  1;
            "HEIGHT_14_59_0": value  <=  2;
            "HEIGHT_14_59_1": value  <=  2;
            "HEIGHT_14_60_0": value  <=  2;
            "HEIGHT_14_60_1": value  <=  2;
            "HEIGHT_14_61_0": value  <=  2;
            "HEIGHT_14_61_1": value  <=  1;
            "HEIGHT_14_62_0": value  <=  4;
            "HEIGHT_14_62_1": value  <=  2;
            "HEIGHT_14_62_2": value  <=  2;
            "HEIGHT_14_63_0": value  <=  3;
            "HEIGHT_14_63_1": value  <=  1;
            "HEIGHT_14_64_0": value  <=  6;
            "HEIGHT_14_64_1": value  <=  2;
            "HEIGHT_14_65_0": value  <=  6;
            "HEIGHT_14_65_1": value  <=  3;
            "HEIGHT_14_66_0": value  <=  3;
            "HEIGHT_14_66_1": value  <=  1;
            "HEIGHT_14_67_0": value  <=  6;
            "HEIGHT_14_67_1": value  <=  2;
            "HEIGHT_14_68_0": value  <=  2;
            "HEIGHT_14_68_1": value  <=  1;
            "HEIGHT_14_69_0": value  <=  2;
            "HEIGHT_14_69_1": value  <=  1;
            "HEIGHT_14_70_0": value  <=  3;
            "HEIGHT_14_70_1": value  <=  1;
            "HEIGHT_14_71_0": value  <=  4;
            "HEIGHT_14_71_1": value  <=  4;
            "HEIGHT_14_72_0": value  <=  1;
            "HEIGHT_14_72_1": value  <=  1;
            "HEIGHT_14_73_0": value  <=  2;
            "HEIGHT_14_73_1": value  <=  2;
            "HEIGHT_14_74_0": value  <=  6;
            "HEIGHT_14_74_1": value  <=  2;
            "HEIGHT_14_75_0": value  <=  3;
            "HEIGHT_14_75_1": value  <=  3;
            "HEIGHT_14_76_0": value  <=  4;
            "HEIGHT_14_76_1": value  <=  4;
            "HEIGHT_14_77_0": value  <=  3;
            "HEIGHT_14_77_1": value  <=  1;
            "HEIGHT_14_78_0": value  <=  2;
            "HEIGHT_14_78_1": value  <=  1;
            "HEIGHT_14_78_2": value  <=  1;
            "HEIGHT_14_79_0": value  <=  5;
            "HEIGHT_14_79_1": value  <=  5;
            "HEIGHT_14_80_0": value  <=  5;
            "HEIGHT_14_80_1": value  <=  5;
            "HEIGHT_14_81_0": value  <=  3;
            "HEIGHT_14_81_1": value  <=  1;
            "HEIGHT_14_82_0": value  <=  3;
            "HEIGHT_14_82_1": value  <=  1;
            "HEIGHT_14_83_0": value  <=  1;
            "HEIGHT_14_83_1": value  <=  1;
            "HEIGHT_14_84_0": value  <=  1;
            "HEIGHT_14_84_1": value  <=  1;
            "HEIGHT_14_85_0": value  <=  3;
            "HEIGHT_14_85_1": value  <=  1;
            "HEIGHT_14_86_0": value  <=  15;
            "HEIGHT_14_86_1": value  <=  15;
            "HEIGHT_14_87_0": value  <=  5;
            "HEIGHT_14_87_1": value  <=  5;
            "HEIGHT_14_88_0": value  <=  7;
            "HEIGHT_14_88_1": value  <=  7;
            "HEIGHT_14_89_0": value  <=  3;
            "HEIGHT_14_89_1": value  <=  1;
            "HEIGHT_14_90_0": value  <=  3;
            "HEIGHT_14_90_1": value  <=  1;
            "HEIGHT_14_91_0": value  <=  3;
            "HEIGHT_14_91_1": value  <=  1;
            "HEIGHT_14_92_0": value  <=  2;
            "HEIGHT_14_92_1": value  <=  1;
            "HEIGHT_14_93_0": value  <=  6;
            "HEIGHT_14_93_1": value  <=  6;
            "HEIGHT_14_94_0": value  <=  4;
            "HEIGHT_14_94_1": value  <=  4;
            "HEIGHT_14_95_0": value  <=  10;
            "HEIGHT_14_95_1": value  <=  5;
            "HEIGHT_14_95_2": value  <=  5;
            "HEIGHT_14_96_0": value  <=  2;
            "HEIGHT_14_96_1": value  <=  2;
            "HEIGHT_14_97_0": value  <=  2;
            "HEIGHT_14_97_1": value  <=  1;
            "HEIGHT_14_98_0": value  <=  10;
            "HEIGHT_14_98_1": value  <=  5;
            "HEIGHT_14_98_2": value  <=  5;
            "HEIGHT_14_99_0": value  <=  6;
            "HEIGHT_14_99_1": value  <=  3;
            "HEIGHT_14_99_2": value  <=  3;
            "HEIGHT_14_100_0": value  <=  15;
            "HEIGHT_14_100_1": value  <=  15;
            "HEIGHT_14_101_0": value  <=  4;
            "HEIGHT_14_101_1": value  <=  2;
            "HEIGHT_14_101_2": value  <=  2;
            "HEIGHT_14_102_0": value  <=  17;
            "HEIGHT_14_102_1": value  <=  17;
            "HEIGHT_14_103_0": value  <=  6;
            "HEIGHT_14_103_1": value  <=  3;
            "HEIGHT_14_103_2": value  <=  3;
            "HEIGHT_14_104_0": value  <=  3;
            "HEIGHT_14_104_1": value  <=  1;
            "HEIGHT_14_105_0": value  <=  2;
            "HEIGHT_14_105_1": value  <=  1;
            "HEIGHT_14_106_0": value  <=  2;
            "HEIGHT_14_106_1": value  <=  1;
            "HEIGHT_14_106_2": value  <=  1;
            "HEIGHT_14_107_0": value  <=  6;
            "HEIGHT_14_107_1": value  <=  3;
            "HEIGHT_14_108_0": value  <=  2;
            "HEIGHT_14_108_1": value  <=  1;
            "HEIGHT_14_109_0": value  <=  6;
            "HEIGHT_14_109_1": value  <=  2;
            "HEIGHT_14_110_0": value  <=  2;
            "HEIGHT_14_110_1": value  <=  1;
            "HEIGHT_14_111_0": value  <=  6;
            "HEIGHT_14_111_1": value  <=  2;
            "HEIGHT_14_112_0": value  <=  3;
            "HEIGHT_14_112_1": value  <=  1;
            "HEIGHT_14_113_0": value  <=  6;
            "HEIGHT_14_113_1": value  <=  2;
            "HEIGHT_14_114_0": value  <=  6;
            "HEIGHT_14_114_1": value  <=  2;
            "HEIGHT_14_115_0": value  <=  3;
            "HEIGHT_14_115_1": value  <=  1;
            "HEIGHT_14_116_0": value  <=  3;
            "HEIGHT_14_116_1": value  <=  1;
            "HEIGHT_14_117_0": value  <=  3;
            "HEIGHT_14_117_1": value  <=  1;
            "HEIGHT_14_118_0": value  <=  3;
            "HEIGHT_14_118_1": value  <=  1;
            "HEIGHT_14_119_0": value  <=  6;
            "HEIGHT_14_119_1": value  <=  2;
            "HEIGHT_14_120_0": value  <=  3;
            "HEIGHT_14_120_1": value  <=  1;
            "HEIGHT_14_121_0": value  <=  5;
            "HEIGHT_14_121_1": value  <=  5;
            "HEIGHT_14_122_0": value  <=  2;
            "HEIGHT_14_122_1": value  <=  2;
            "HEIGHT_14_123_0": value  <=  9;
            "HEIGHT_14_123_1": value  <=  9;
            "HEIGHT_14_124_0": value  <=  6;
            "HEIGHT_14_124_1": value  <=  6;
            "HEIGHT_14_125_0": value  <=  3;
            "HEIGHT_14_125_1": value  <=  1;
            "HEIGHT_14_126_0": value  <=  9;
            "HEIGHT_14_126_1": value  <=  9;
            "HEIGHT_14_127_0": value  <=  5;
            "HEIGHT_14_127_1": value  <=  5;
            "HEIGHT_14_128_0": value  <=  3;
            "HEIGHT_14_128_1": value  <=  3;
            "HEIGHT_14_129_0": value  <=  5;
            "HEIGHT_14_129_1": value  <=  5;
            "HEIGHT_14_130_0": value  <=  2;
            "HEIGHT_14_130_1": value  <=  2;
            "HEIGHT_14_131_0": value  <=  2;
            "HEIGHT_14_131_1": value  <=  2;
            "HEIGHT_14_132_0": value  <=  3;
            "HEIGHT_14_132_1": value  <=  3;
            "HEIGHT_14_133_0": value  <=  1;
            "HEIGHT_14_133_1": value  <=  1;
            "HEIGHT_14_134_0": value  <=  15;
            "HEIGHT_14_134_1": value  <=  5;
            "HEIGHT_15_0_0": value  <=  6;
            "HEIGHT_15_0_1": value  <=  6;
            "HEIGHT_15_1_0": value  <=  1;
            "HEIGHT_15_1_1": value  <=  1;
            "HEIGHT_15_2_0": value  <=  4;
            "HEIGHT_15_2_1": value  <=  2;
            "HEIGHT_15_2_2": value  <=  2;
            "HEIGHT_15_3_0": value  <=  8;
            "HEIGHT_15_3_1": value  <=  4;
            "HEIGHT_15_4_0": value  <=  6;
            "HEIGHT_15_4_1": value  <=  3;
            "HEIGHT_15_5_0": value  <=  10;
            "HEIGHT_15_5_1": value  <=  5;
            "HEIGHT_15_5_2": value  <=  5;
            "HEIGHT_15_6_0": value  <=  10;
            "HEIGHT_15_6_1": value  <=  5;
            "HEIGHT_15_6_2": value  <=  5;
            "HEIGHT_15_7_0": value  <=  2;
            "HEIGHT_15_7_1": value  <=  1;
            "HEIGHT_15_8_0": value  <=  2;
            "HEIGHT_15_8_1": value  <=  1;
            "HEIGHT_15_9_0": value  <=  2;
            "HEIGHT_15_9_1": value  <=  1;
            "HEIGHT_15_10_0": value  <=  10;
            "HEIGHT_15_10_1": value  <=  5;
            "HEIGHT_15_10_2": value  <=  5;
            "HEIGHT_15_11_0": value  <=  2;
            "HEIGHT_15_11_1": value  <=  1;
            "HEIGHT_15_12_0": value  <=  3;
            "HEIGHT_15_12_1": value  <=  1;
            "HEIGHT_15_13_0": value  <=  3;
            "HEIGHT_15_13_1": value  <=  1;
            "HEIGHT_15_14_0": value  <=  2;
            "HEIGHT_15_14_1": value  <=  2;
            "HEIGHT_15_15_0": value  <=  3;
            "HEIGHT_15_15_1": value  <=  1;
            "HEIGHT_15_16_0": value  <=  2;
            "HEIGHT_15_16_1": value  <=  1;
            "HEIGHT_15_17_0": value  <=  6;
            "HEIGHT_15_17_1": value  <=  2;
            "HEIGHT_15_18_0": value  <=  4;
            "HEIGHT_15_18_1": value  <=  4;
            "HEIGHT_15_19_0": value  <=  6;
            "HEIGHT_15_19_1": value  <=  2;
            "HEIGHT_15_20_0": value  <=  8;
            "HEIGHT_15_20_1": value  <=  8;
            "HEIGHT_15_21_0": value  <=  6;
            "HEIGHT_15_21_1": value  <=  3;
            "HEIGHT_15_22_0": value  <=  2;
            "HEIGHT_15_22_1": value  <=  1;
            "HEIGHT_15_23_0": value  <=  6;
            "HEIGHT_15_23_1": value  <=  2;
            "HEIGHT_15_24_0": value  <=  6;
            "HEIGHT_15_24_1": value  <=  2;
            "HEIGHT_15_25_0": value  <=  6;
            "HEIGHT_15_25_1": value  <=  3;
            "HEIGHT_15_26_0": value  <=  6;
            "HEIGHT_15_26_1": value  <=  6;
            "HEIGHT_15_27_0": value  <=  6;
            "HEIGHT_15_27_1": value  <=  3;
            "HEIGHT_15_27_2": value  <=  3;
            "HEIGHT_15_28_0": value  <=  5;
            "HEIGHT_15_28_1": value  <=  5;
            "HEIGHT_15_29_0": value  <=  6;
            "HEIGHT_15_29_1": value  <=  2;
            "HEIGHT_15_30_0": value  <=  5;
            "HEIGHT_15_30_1": value  <=  5;
            "HEIGHT_15_31_0": value  <=  2;
            "HEIGHT_15_31_1": value  <=  2;
            "HEIGHT_15_32_0": value  <=  2;
            "HEIGHT_15_32_1": value  <=  2;
            "HEIGHT_15_33_0": value  <=  2;
            "HEIGHT_15_33_1": value  <=  1;
            "HEIGHT_15_34_0": value  <=  12;
            "HEIGHT_15_34_1": value  <=  6;
            "HEIGHT_15_35_0": value  <=  4;
            "HEIGHT_15_35_1": value  <=  4;
            "HEIGHT_15_36_0": value  <=  2;
            "HEIGHT_15_36_1": value  <=  1;
            "HEIGHT_15_37_0": value  <=  2;
            "HEIGHT_15_37_1": value  <=  1;
            "HEIGHT_15_37_2": value  <=  1;
            "HEIGHT_15_38_0": value  <=  6;
            "HEIGHT_15_38_1": value  <=  2;
            "HEIGHT_15_39_0": value  <=  3;
            "HEIGHT_15_39_1": value  <=  1;
            "HEIGHT_15_40_0": value  <=  3;
            "HEIGHT_15_40_1": value  <=  1;
            "HEIGHT_15_41_0": value  <=  1;
            "HEIGHT_15_41_1": value  <=  1;
            "HEIGHT_15_42_0": value  <=  1;
            "HEIGHT_15_42_1": value  <=  1;
            "HEIGHT_15_43_0": value  <=  3;
            "HEIGHT_15_43_1": value  <=  1;
            "HEIGHT_15_44_0": value  <=  3;
            "HEIGHT_15_44_1": value  <=  1;
            "HEIGHT_15_45_0": value  <=  3;
            "HEIGHT_15_45_1": value  <=  1;
            "HEIGHT_15_46_0": value  <=  3;
            "HEIGHT_15_46_1": value  <=  1;
            "HEIGHT_15_47_0": value  <=  3;
            "HEIGHT_15_47_1": value  <=  1;
            "HEIGHT_15_48_0": value  <=  3;
            "HEIGHT_15_48_1": value  <=  3;
            "HEIGHT_15_49_0": value  <=  17;
            "HEIGHT_15_49_1": value  <=  17;
            "HEIGHT_15_50_0": value  <=  3;
            "HEIGHT_15_50_1": value  <=  1;
            "HEIGHT_15_51_0": value  <=  15;
            "HEIGHT_15_51_1": value  <=  5;
            "HEIGHT_15_52_0": value  <=  3;
            "HEIGHT_15_52_1": value  <=  1;
            "HEIGHT_15_53_0": value  <=  3;
            "HEIGHT_15_53_1": value  <=  1;
            "HEIGHT_15_54_0": value  <=  5;
            "HEIGHT_15_54_1": value  <=  5;
            "HEIGHT_15_55_0": value  <=  2;
            "HEIGHT_15_55_1": value  <=  2;
            "HEIGHT_15_56_0": value  <=  3;
            "HEIGHT_15_56_1": value  <=  1;
            "HEIGHT_15_57_0": value  <=  3;
            "HEIGHT_15_57_1": value  <=  1;
            "HEIGHT_15_58_0": value  <=  15;
            "HEIGHT_15_58_1": value  <=  5;
            "HEIGHT_15_59_0": value  <=  10;
            "HEIGHT_15_59_1": value  <=  5;
            "HEIGHT_15_59_2": value  <=  5;
            "HEIGHT_15_60_0": value  <=  3;
            "HEIGHT_15_60_1": value  <=  3;
            "HEIGHT_15_61_0": value  <=  1;
            "HEIGHT_15_61_1": value  <=  1;
            "HEIGHT_15_62_0": value  <=  10;
            "HEIGHT_15_62_1": value  <=  5;
            "HEIGHT_15_62_2": value  <=  5;
            "HEIGHT_15_63_0": value  <=  1;
            "HEIGHT_15_63_1": value  <=  1;
            "HEIGHT_15_64_0": value  <=  6;
            "HEIGHT_15_64_1": value  <=  2;
            "HEIGHT_15_65_0": value  <=  1;
            "HEIGHT_15_65_1": value  <=  1;
            "HEIGHT_15_66_0": value  <=  1;
            "HEIGHT_15_66_1": value  <=  1;
            "HEIGHT_15_67_0": value  <=  4;
            "HEIGHT_15_67_1": value  <=  2;
            "HEIGHT_15_67_2": value  <=  2;
            "HEIGHT_15_68_0": value  <=  2;
            "HEIGHT_15_68_1": value  <=  1;
            "HEIGHT_15_68_2": value  <=  1;
            "HEIGHT_15_69_0": value  <=  2;
            "HEIGHT_15_69_1": value  <=  1;
            "HEIGHT_15_70_0": value  <=  18;
            "HEIGHT_15_70_1": value  <=  9;
            "HEIGHT_15_70_2": value  <=  9;
            "HEIGHT_15_71_0": value  <=  4;
            "HEIGHT_15_71_1": value  <=  2;
            "HEIGHT_15_71_2": value  <=  2;
            "HEIGHT_15_72_0": value  <=  3;
            "HEIGHT_15_72_1": value  <=  1;
            "HEIGHT_15_73_0": value  <=  4;
            "HEIGHT_15_73_1": value  <=  2;
            "HEIGHT_15_73_2": value  <=  2;
            "HEIGHT_15_74_0": value  <=  4;
            "HEIGHT_15_74_1": value  <=  2;
            "HEIGHT_15_74_2": value  <=  2;
            "HEIGHT_15_75_0": value  <=  3;
            "HEIGHT_15_75_1": value  <=  1;
            "HEIGHT_15_76_0": value  <=  3;
            "HEIGHT_15_76_1": value  <=  1;
            "HEIGHT_15_77_0": value  <=  3;
            "HEIGHT_15_77_1": value  <=  1;
            "HEIGHT_15_78_0": value  <=  4;
            "HEIGHT_15_78_1": value  <=  4;
            "HEIGHT_15_79_0": value  <=  4;
            "HEIGHT_15_79_1": value  <=  4;
            "HEIGHT_15_80_0": value  <=  3;
            "HEIGHT_15_80_1": value  <=  3;
            "HEIGHT_15_81_0": value  <=  8;
            "HEIGHT_15_81_1": value  <=  4;
            "HEIGHT_15_81_2": value  <=  4;
            "HEIGHT_15_82_0": value  <=  12;
            "HEIGHT_15_82_1": value  <=  6;
            "HEIGHT_15_82_2": value  <=  6;
            "HEIGHT_15_83_0": value  <=  12;
            "HEIGHT_15_83_1": value  <=  6;
            "HEIGHT_15_84_0": value  <=  14;
            "HEIGHT_15_84_1": value  <=  7;
            "HEIGHT_15_85_0": value  <=  1;
            "HEIGHT_15_85_1": value  <=  1;
            "HEIGHT_15_86_0": value  <=  4;
            "HEIGHT_15_86_1": value  <=  2;
            "HEIGHT_15_87_0": value  <=  8;
            "HEIGHT_15_87_1": value  <=  4;
            "HEIGHT_15_88_0": value  <=  8;
            "HEIGHT_15_88_1": value  <=  4;
            "HEIGHT_15_88_2": value  <=  4;
            "HEIGHT_15_89_0": value  <=  1;
            "HEIGHT_15_89_1": value  <=  1;
            "HEIGHT_15_90_0": value  <=  4;
            "HEIGHT_15_90_1": value  <=  4;
            "HEIGHT_15_91_0": value  <=  6;
            "HEIGHT_15_91_1": value  <=  2;
            "HEIGHT_15_92_0": value  <=  4;
            "HEIGHT_15_92_1": value  <=  4;
            "HEIGHT_15_93_0": value  <=  3;
            "HEIGHT_15_93_1": value  <=  1;
            "HEIGHT_15_94_0": value  <=  1;
            "HEIGHT_15_94_1": value  <=  1;
            "HEIGHT_15_95_0": value  <=  6;
            "HEIGHT_15_95_1": value  <=  2;
            "HEIGHT_15_96_0": value  <=  1;
            "HEIGHT_15_96_1": value  <=  1;
            "HEIGHT_15_97_0": value  <=  10;
            "HEIGHT_15_97_1": value  <=  5;
            "HEIGHT_15_97_2": value  <=  5;
            "HEIGHT_15_98_0": value  <=  9;
            "HEIGHT_15_98_1": value  <=  3;
            "HEIGHT_15_99_0": value  <=  3;
            "HEIGHT_15_99_1": value  <=  1;
            "HEIGHT_15_100_0": value  <=  3;
            "HEIGHT_15_100_1": value  <=  3;
            "HEIGHT_15_101_0": value  <=  3;
            "HEIGHT_15_101_1": value  <=  1;
            "HEIGHT_15_102_0": value  <=  10;
            "HEIGHT_15_102_1": value  <=  10;
            "HEIGHT_15_103_0": value  <=  3;
            "HEIGHT_15_103_1": value  <=  1;
            "HEIGHT_15_104_0": value  <=  6;
            "HEIGHT_15_104_1": value  <=  2;
            "HEIGHT_15_105_0": value  <=  3;
            "HEIGHT_15_105_1": value  <=  1;
            "HEIGHT_15_106_0": value  <=  3;
            "HEIGHT_15_106_1": value  <=  1;
            "HEIGHT_15_107_0": value  <=  8;
            "HEIGHT_15_107_1": value  <=  4;
            "HEIGHT_15_107_2": value  <=  4;
            "HEIGHT_15_108_0": value  <=  8;
            "HEIGHT_15_108_1": value  <=  4;
            "HEIGHT_15_108_2": value  <=  4;
            "HEIGHT_15_109_0": value  <=  10;
            "HEIGHT_15_109_1": value  <=  5;
            "HEIGHT_15_109_2": value  <=  5;
            "HEIGHT_15_110_0": value  <=  3;
            "HEIGHT_15_110_1": value  <=  1;
            "HEIGHT_15_111_0": value  <=  3;
            "HEIGHT_15_111_1": value  <=  1;
            "HEIGHT_15_112_0": value  <=  3;
            "HEIGHT_15_112_1": value  <=  1;
            "HEIGHT_15_113_0": value  <=  3;
            "HEIGHT_15_113_1": value  <=  1;
            "HEIGHT_15_114_0": value  <=  3;
            "HEIGHT_15_114_1": value  <=  1;
            "HEIGHT_15_115_0": value  <=  2;
            "HEIGHT_15_115_1": value  <=  1;
            "HEIGHT_15_116_0": value  <=  12;
            "HEIGHT_15_116_1": value  <=  12;
            "HEIGHT_15_117_0": value  <=  3;
            "HEIGHT_15_117_1": value  <=  1;
            "HEIGHT_15_118_0": value  <=  4;
            "HEIGHT_15_118_1": value  <=  2;
            "HEIGHT_15_119_0": value  <=  14;
            "HEIGHT_15_119_1": value  <=  7;
            "HEIGHT_15_120_0": value  <=  10;
            "HEIGHT_15_120_1": value  <=  5;
            "HEIGHT_15_120_2": value  <=  5;
            "HEIGHT_15_121_0": value  <=  4;
            "HEIGHT_15_121_1": value  <=  4;
            "HEIGHT_15_122_0": value  <=  4;
            "HEIGHT_15_122_1": value  <=  4;
            "HEIGHT_15_123_0": value  <=  2;
            "HEIGHT_15_123_1": value  <=  1;
            "HEIGHT_15_124_0": value  <=  2;
            "HEIGHT_15_124_1": value  <=  1;
            "HEIGHT_15_125_0": value  <=  2;
            "HEIGHT_15_125_1": value  <=  1;
            "HEIGHT_15_125_2": value  <=  1;
            "HEIGHT_15_126_0": value  <=  2;
            "HEIGHT_15_126_1": value  <=  1;
            "HEIGHT_15_126_2": value  <=  1;
            "HEIGHT_15_127_0": value  <=  3;
            "HEIGHT_15_127_1": value  <=  3;
            "HEIGHT_15_128_0": value  <=  12;
            "HEIGHT_15_128_1": value  <=  12;
            "HEIGHT_15_129_0": value  <=  3;
            "HEIGHT_15_129_1": value  <=  1;
            "HEIGHT_15_130_0": value  <=  3;
            "HEIGHT_15_130_1": value  <=  1;
            "HEIGHT_15_131_0": value  <=  3;
            "HEIGHT_15_131_1": value  <=  1;
            "HEIGHT_15_132_0": value  <=  3;
            "HEIGHT_15_132_1": value  <=  1;
            "HEIGHT_15_133_0": value  <=  6;
            "HEIGHT_15_133_1": value  <=  3;
            "HEIGHT_15_133_2": value  <=  3;
            "HEIGHT_15_134_0": value  <=  3;
            "HEIGHT_15_134_1": value  <=  1;
            "HEIGHT_15_135_0": value  <=  20;
            "HEIGHT_15_135_1": value  <=  20;
            "HEIGHT_15_136_0": value  <=  6;
            "HEIGHT_15_136_1": value  <=  3;
            "HEIGHT_15_136_2": value  <=  3;
            "HEIGHT_16_0_0": value  <=  4;
            "HEIGHT_16_0_1": value  <=  2;
            "HEIGHT_16_1_0": value  <=  12;
            "HEIGHT_16_1_1": value  <=  12;
            "HEIGHT_16_2_0": value  <=  12;
            "HEIGHT_16_2_1": value  <=  6;
            "HEIGHT_16_3_0": value  <=  8;
            "HEIGHT_16_3_1": value  <=  4;
            "HEIGHT_16_4_0": value  <=  10;
            "HEIGHT_16_4_1": value  <=  5;
            "HEIGHT_16_4_2": value  <=  5;
            "HEIGHT_16_5_0": value  <=  14;
            "HEIGHT_16_5_1": value  <=  7;
            "HEIGHT_16_5_2": value  <=  7;
            "HEIGHT_16_6_0": value  <=  14;
            "HEIGHT_16_6_1": value  <=  7;
            "HEIGHT_16_6_2": value  <=  7;
            "HEIGHT_16_7_0": value  <=  2;
            "HEIGHT_16_7_1": value  <=  2;
            "HEIGHT_16_8_0": value  <=  3;
            "HEIGHT_16_8_1": value  <=  1;
            "HEIGHT_16_9_0": value  <=  4;
            "HEIGHT_16_9_1": value  <=  2;
            "HEIGHT_16_9_2": value  <=  2;
            "HEIGHT_16_10_0": value  <=  2;
            "HEIGHT_16_10_1": value  <=  2;
            "HEIGHT_16_11_0": value  <=  9;
            "HEIGHT_16_11_1": value  <=  3;
            "HEIGHT_16_12_0": value  <=  8;
            "HEIGHT_16_12_1": value  <=  8;
            "HEIGHT_16_13_0": value  <=  6;
            "HEIGHT_16_13_1": value  <=  3;
            "HEIGHT_16_14_0": value  <=  4;
            "HEIGHT_16_14_1": value  <=  2;
            "HEIGHT_16_14_2": value  <=  2;
            "HEIGHT_16_15_0": value  <=  19;
            "HEIGHT_16_15_1": value  <=  19;
            "HEIGHT_16_16_0": value  <=  5;
            "HEIGHT_16_16_1": value  <=  5;
            "HEIGHT_16_17_0": value  <=  2;
            "HEIGHT_16_17_1": value  <=  1;
            "HEIGHT_16_18_0": value  <=  2;
            "HEIGHT_16_18_1": value  <=  1;
            "HEIGHT_16_19_0": value  <=  6;
            "HEIGHT_16_19_1": value  <=  2;
            "HEIGHT_16_20_0": value  <=  3;
            "HEIGHT_16_20_1": value  <=  1;
            "HEIGHT_16_21_0": value  <=  6;
            "HEIGHT_16_21_1": value  <=  3;
            "HEIGHT_16_22_0": value  <=  3;
            "HEIGHT_16_22_1": value  <=  1;
            "HEIGHT_16_23_0": value  <=  6;
            "HEIGHT_16_23_1": value  <=  2;
            "HEIGHT_16_24_0": value  <=  3;
            "HEIGHT_16_24_1": value  <=  1;
            "HEIGHT_16_25_0": value  <=  2;
            "HEIGHT_16_25_1": value  <=  2;
            "HEIGHT_16_26_0": value  <=  6;
            "HEIGHT_16_26_1": value  <=  2;
            "HEIGHT_16_27_0": value  <=  6;
            "HEIGHT_16_27_1": value  <=  2;
            "HEIGHT_16_28_0": value  <=  2;
            "HEIGHT_16_28_1": value  <=  1;
            "HEIGHT_16_29_0": value  <=  4;
            "HEIGHT_16_29_1": value  <=  4;
            "HEIGHT_16_30_0": value  <=  9;
            "HEIGHT_16_30_1": value  <=  3;
            "HEIGHT_16_31_0": value  <=  3;
            "HEIGHT_16_31_1": value  <=  1;
            "HEIGHT_16_32_0": value  <=  3;
            "HEIGHT_16_32_1": value  <=  3;
            "HEIGHT_16_33_0": value  <=  8;
            "HEIGHT_16_33_1": value  <=  4;
            "HEIGHT_16_34_0": value  <=  3;
            "HEIGHT_16_34_1": value  <=  1;
            "HEIGHT_16_35_0": value  <=  2;
            "HEIGHT_16_35_1": value  <=  1;
            "HEIGHT_16_35_2": value  <=  1;
            "HEIGHT_16_36_0": value  <=  2;
            "HEIGHT_16_36_1": value  <=  1;
            "HEIGHT_16_36_2": value  <=  1;
            "HEIGHT_16_37_0": value  <=  4;
            "HEIGHT_16_37_1": value  <=  4;
            "HEIGHT_16_38_0": value  <=  7;
            "HEIGHT_16_38_1": value  <=  7;
            "HEIGHT_16_39_0": value  <=  14;
            "HEIGHT_16_39_1": value  <=  7;
            "HEIGHT_16_40_0": value  <=  2;
            "HEIGHT_16_40_1": value  <=  2;
            "HEIGHT_16_41_0": value  <=  4;
            "HEIGHT_16_41_1": value  <=  2;
            "HEIGHT_16_41_2": value  <=  2;
            "HEIGHT_16_42_0": value  <=  2;
            "HEIGHT_16_42_1": value  <=  2;
            "HEIGHT_16_43_0": value  <=  3;
            "HEIGHT_16_43_1": value  <=  3;
            "HEIGHT_16_44_0": value  <=  2;
            "HEIGHT_16_44_1": value  <=  2;
            "HEIGHT_16_45_0": value  <=  7;
            "HEIGHT_16_45_1": value  <=  7;
            "HEIGHT_16_46_0": value  <=  3;
            "HEIGHT_16_46_1": value  <=  3;
            "HEIGHT_16_47_0": value  <=  18;
            "HEIGHT_16_47_1": value  <=  9;
            "HEIGHT_16_48_0": value  <=  3;
            "HEIGHT_16_48_1": value  <=  1;
            "HEIGHT_16_49_0": value  <=  6;
            "HEIGHT_16_49_1": value  <=  6;
            "HEIGHT_16_50_0": value  <=  3;
            "HEIGHT_16_50_1": value  <=  1;
            "HEIGHT_16_51_0": value  <=  3;
            "HEIGHT_16_51_1": value  <=  1;
            "HEIGHT_16_52_0": value  <=  3;
            "HEIGHT_16_52_1": value  <=  1;
            "HEIGHT_16_53_0": value  <=  2;
            "HEIGHT_16_53_1": value  <=  2;
            "HEIGHT_16_54_0": value  <=  6;
            "HEIGHT_16_54_1": value  <=  3;
            "HEIGHT_16_55_0": value  <=  2;
            "HEIGHT_16_55_1": value  <=  1;
            "HEIGHT_16_56_0": value  <=  6;
            "HEIGHT_16_56_1": value  <=  3;
            "HEIGHT_16_56_2": value  <=  3;
            "HEIGHT_16_57_0": value  <=  4;
            "HEIGHT_16_57_1": value  <=  2;
            "HEIGHT_16_58_0": value  <=  3;
            "HEIGHT_16_58_1": value  <=  1;
            "HEIGHT_16_59_0": value  <=  9;
            "HEIGHT_16_59_1": value  <=  3;
            "HEIGHT_16_60_0": value  <=  6;
            "HEIGHT_16_60_1": value  <=  2;
            "HEIGHT_16_61_0": value  <=  6;
            "HEIGHT_16_61_1": value  <=  3;
            "HEIGHT_16_62_0": value  <=  8;
            "HEIGHT_16_62_1": value  <=  8;
            "HEIGHT_16_63_0": value  <=  18;
            "HEIGHT_16_63_1": value  <=  18;
            "HEIGHT_16_64_0": value  <=  2;
            "HEIGHT_16_64_1": value  <=  1;
            "HEIGHT_16_65_0": value  <=  6;
            "HEIGHT_16_65_1": value  <=  2;
            "HEIGHT_16_66_0": value  <=  6;
            "HEIGHT_16_66_1": value  <=  3;
            "HEIGHT_16_67_0": value  <=  3;
            "HEIGHT_16_67_1": value  <=  1;
            "HEIGHT_16_68_0": value  <=  18;
            "HEIGHT_16_68_1": value  <=  18;
            "HEIGHT_16_69_0": value  <=  2;
            "HEIGHT_16_69_1": value  <=  1;
            "HEIGHT_16_69_2": value  <=  1;
            "HEIGHT_16_70_0": value  <=  2;
            "HEIGHT_16_70_1": value  <=  1;
            "HEIGHT_16_71_0": value  <=  3;
            "HEIGHT_16_71_1": value  <=  1;
            "HEIGHT_16_72_0": value  <=  3;
            "HEIGHT_16_72_1": value  <=  1;
            "HEIGHT_16_73_0": value  <=  3;
            "HEIGHT_16_73_1": value  <=  3;
            "HEIGHT_16_74_0": value  <=  2;
            "HEIGHT_16_74_1": value  <=  2;
            "HEIGHT_16_75_0": value  <=  2;
            "HEIGHT_16_75_1": value  <=  1;
            "HEIGHT_16_76_0": value  <=  2;
            "HEIGHT_16_76_1": value  <=  1;
            "HEIGHT_16_77_0": value  <=  6;
            "HEIGHT_16_77_1": value  <=  3;
            "HEIGHT_16_78_0": value  <=  3;
            "HEIGHT_16_78_1": value  <=  3;
            "HEIGHT_16_79_0": value  <=  3;
            "HEIGHT_16_79_1": value  <=  3;
            "HEIGHT_16_80_0": value  <=  18;
            "HEIGHT_16_80_1": value  <=  18;
            "HEIGHT_16_81_0": value  <=  3;
            "HEIGHT_16_81_1": value  <=  1;
            "HEIGHT_16_82_0": value  <=  6;
            "HEIGHT_16_82_1": value  <=  3;
            "HEIGHT_16_83_0": value  <=  2;
            "HEIGHT_16_83_1": value  <=  1;
            "HEIGHT_16_84_0": value  <=  3;
            "HEIGHT_16_84_1": value  <=  3;
            "HEIGHT_16_85_0": value  <=  3;
            "HEIGHT_16_85_1": value  <=  1;
            "HEIGHT_16_86_0": value  <=  3;
            "HEIGHT_16_86_1": value  <=  1;
            "HEIGHT_16_87_0": value  <=  2;
            "HEIGHT_16_87_1": value  <=  1;
            "HEIGHT_16_87_2": value  <=  1;
            "HEIGHT_16_88_0": value  <=  2;
            "HEIGHT_16_88_1": value  <=  1;
            "HEIGHT_16_88_2": value  <=  1;
            "HEIGHT_16_89_0": value  <=  4;
            "HEIGHT_16_89_1": value  <=  2;
            "HEIGHT_16_90_0": value  <=  4;
            "HEIGHT_16_90_1": value  <=  2;
            "HEIGHT_16_91_0": value  <=  3;
            "HEIGHT_16_91_1": value  <=  1;
            "HEIGHT_16_92_0": value  <=  20;
            "HEIGHT_16_92_1": value  <=  20;
            "HEIGHT_16_93_0": value  <=  8;
            "HEIGHT_16_93_1": value  <=  4;
            "HEIGHT_16_93_2": value  <=  4;
            "HEIGHT_16_94_0": value  <=  2;
            "HEIGHT_16_94_1": value  <=  1;
            "HEIGHT_16_94_2": value  <=  1;
            "HEIGHT_16_95_0": value  <=  3;
            "HEIGHT_16_95_1": value  <=  1;
            "HEIGHT_16_96_0": value  <=  2;
            "HEIGHT_16_96_1": value  <=  1;
            "HEIGHT_16_97_0": value  <=  12;
            "HEIGHT_16_97_1": value  <=  6;
            "HEIGHT_16_98_0": value  <=  12;
            "HEIGHT_16_98_1": value  <=  4;
            "HEIGHT_16_99_0": value  <=  11;
            "HEIGHT_16_99_1": value  <=  11;
            "HEIGHT_16_100_0": value  <=  3;
            "HEIGHT_16_100_1": value  <=  1;
            "HEIGHT_16_101_0": value  <=  3;
            "HEIGHT_16_101_1": value  <=  1;
            "HEIGHT_16_102_0": value  <=  2;
            "HEIGHT_16_102_1": value  <=  1;
            "HEIGHT_16_103_0": value  <=  3;
            "HEIGHT_16_103_1": value  <=  3;
            "HEIGHT_16_104_0": value  <=  4;
            "HEIGHT_16_104_1": value  <=  4;
            "HEIGHT_16_105_0": value  <=  3;
            "HEIGHT_16_105_1": value  <=  3;
            "HEIGHT_16_106_0": value  <=  2;
            "HEIGHT_16_106_1": value  <=  2;
            "HEIGHT_16_107_0": value  <=  4;
            "HEIGHT_16_107_1": value  <=  2;
            "HEIGHT_16_107_2": value  <=  2;
            "HEIGHT_16_108_0": value  <=  17;
            "HEIGHT_16_108_1": value  <=  17;
            "HEIGHT_16_109_0": value  <=  7;
            "HEIGHT_16_109_1": value  <=  7;
            "HEIGHT_16_110_0": value  <=  1;
            "HEIGHT_16_110_1": value  <=  1;
            "HEIGHT_16_111_0": value  <=  4;
            "HEIGHT_16_111_1": value  <=  4;
            "HEIGHT_16_112_0": value  <=  12;
            "HEIGHT_16_112_1": value  <=  6;
            "HEIGHT_16_112_2": value  <=  6;
            "HEIGHT_16_113_0": value  <=  2;
            "HEIGHT_16_113_1": value  <=  1;
            "HEIGHT_16_113_2": value  <=  1;
            "HEIGHT_16_114_0": value  <=  6;
            "HEIGHT_16_114_1": value  <=  2;
            "HEIGHT_16_115_0": value  <=  3;
            "HEIGHT_16_115_1": value  <=  3;
            "HEIGHT_16_116_0": value  <=  12;
            "HEIGHT_16_116_1": value  <=  12;
            "HEIGHT_16_117_0": value  <=  2;
            "HEIGHT_16_117_1": value  <=  2;
            "HEIGHT_16_118_0": value  <=  3;
            "HEIGHT_16_118_1": value  <=  1;
            "HEIGHT_16_119_0": value  <=  3;
            "HEIGHT_16_119_1": value  <=  1;
            "HEIGHT_16_120_0": value  <=  6;
            "HEIGHT_16_120_1": value  <=  2;
            "HEIGHT_16_121_0": value  <=  3;
            "HEIGHT_16_121_1": value  <=  1;
            "HEIGHT_16_122_0": value  <=  3;
            "HEIGHT_16_122_1": value  <=  1;
            "HEIGHT_16_123_0": value  <=  1;
            "HEIGHT_16_123_1": value  <=  1;
            "HEIGHT_16_124_0": value  <=  19;
            "HEIGHT_16_124_1": value  <=  19;
            "HEIGHT_16_125_0": value  <=  6;
            "HEIGHT_16_125_1": value  <=  3;
            "HEIGHT_16_125_2": value  <=  3;
            "HEIGHT_16_126_0": value  <=  2;
            "HEIGHT_16_126_1": value  <=  1;
            "HEIGHT_16_126_2": value  <=  1;
            "HEIGHT_16_127_0": value  <=  2;
            "HEIGHT_16_127_1": value  <=  1;
            "HEIGHT_16_127_2": value  <=  1;
            "HEIGHT_16_128_0": value  <=  2;
            "HEIGHT_16_128_1": value  <=  1;
            "HEIGHT_16_128_2": value  <=  1;
            "HEIGHT_16_129_0": value  <=  12;
            "HEIGHT_16_129_1": value  <=  6;
            "HEIGHT_16_130_0": value  <=  10;
            "HEIGHT_16_130_1": value  <=  5;
            "HEIGHT_16_130_2": value  <=  5;
            "HEIGHT_16_131_0": value  <=  2;
            "HEIGHT_16_131_1": value  <=  2;
            "HEIGHT_16_132_0": value  <=  2;
            "HEIGHT_16_132_1": value  <=  1;
            "HEIGHT_16_133_0": value  <=  5;
            "HEIGHT_16_133_1": value  <=  5;
            "HEIGHT_16_134_0": value  <=  5;
            "HEIGHT_16_134_1": value  <=  5;
            "HEIGHT_16_135_0": value  <=  17;
            "HEIGHT_16_135_1": value  <=  17;
            "HEIGHT_16_136_0": value  <=  17;
            "HEIGHT_16_136_1": value  <=  17;
            "HEIGHT_16_137_0": value  <=  9;
            "HEIGHT_16_137_1": value  <=  9;
            "HEIGHT_16_138_0": value  <=  9;
            "HEIGHT_16_138_1": value  <=  9;
            "HEIGHT_16_139_0": value  <=  4;
            "HEIGHT_16_139_1": value  <=  4;
            "HEIGHT_17_0_0": value  <=  1;
            "HEIGHT_17_0_1": value  <=  1;
            "HEIGHT_17_1_0": value  <=  4;
            "HEIGHT_17_1_1": value  <=  2;
            "HEIGHT_17_1_2": value  <=  2;
            "HEIGHT_17_2_0": value  <=  12;
            "HEIGHT_17_2_1": value  <=  4;
            "HEIGHT_17_3_0": value  <=  6;
            "HEIGHT_17_3_1": value  <=  2;
            "HEIGHT_17_4_0": value  <=  6;
            "HEIGHT_17_4_1": value  <=  3;
            "HEIGHT_17_4_2": value  <=  3;
            "HEIGHT_17_5_0": value  <=  4;
            "HEIGHT_17_5_1": value  <=  2;
            "HEIGHT_17_5_2": value  <=  2;
            "HEIGHT_17_6_0": value  <=  3;
            "HEIGHT_17_6_1": value  <=  3;
            "HEIGHT_17_7_0": value  <=  10;
            "HEIGHT_17_7_1": value  <=  5;
            "HEIGHT_17_8_0": value  <=  4;
            "HEIGHT_17_8_1": value  <=  4;
            "HEIGHT_17_9_0": value  <=  6;
            "HEIGHT_17_9_1": value  <=  3;
            "HEIGHT_17_10_0": value  <=  3;
            "HEIGHT_17_10_1": value  <=  1;
            "HEIGHT_17_11_0": value  <=  6;
            "HEIGHT_17_11_1": value  <=  3;
            "HEIGHT_17_11_2": value  <=  3;
            "HEIGHT_17_12_0": value  <=  9;
            "HEIGHT_17_12_1": value  <=  3;
            "HEIGHT_17_13_0": value  <=  6;
            "HEIGHT_17_13_1": value  <=  2;
            "HEIGHT_17_14_0": value  <=  6;
            "HEIGHT_17_14_1": value  <=  2;
            "HEIGHT_17_15_0": value  <=  3;
            "HEIGHT_17_15_1": value  <=  1;
            "HEIGHT_17_16_0": value  <=  6;
            "HEIGHT_17_16_1": value  <=  2;
            "HEIGHT_17_17_0": value  <=  3;
            "HEIGHT_17_17_1": value  <=  1;
            "HEIGHT_17_18_0": value  <=  3;
            "HEIGHT_17_18_1": value  <=  3;
            "HEIGHT_17_19_0": value  <=  3;
            "HEIGHT_17_19_1": value  <=  1;
            "HEIGHT_17_20_0": value  <=  3;
            "HEIGHT_17_20_1": value  <=  1;
            "HEIGHT_17_21_0": value  <=  2;
            "HEIGHT_17_21_1": value  <=  1;
            "HEIGHT_17_22_0": value  <=  6;
            "HEIGHT_17_22_1": value  <=  6;
            "HEIGHT_17_23_0": value  <=  1;
            "HEIGHT_17_23_1": value  <=  1;
            "HEIGHT_17_24_0": value  <=  1;
            "HEIGHT_17_24_1": value  <=  1;
            "HEIGHT_17_25_0": value  <=  5;
            "HEIGHT_17_25_1": value  <=  5;
            "HEIGHT_17_26_0": value  <=  2;
            "HEIGHT_17_26_1": value  <=  2;
            "HEIGHT_17_27_0": value  <=  3;
            "HEIGHT_17_27_1": value  <=  1;
            "HEIGHT_17_28_0": value  <=  1;
            "HEIGHT_17_28_1": value  <=  1;
            "HEIGHT_17_29_0": value  <=  3;
            "HEIGHT_17_29_1": value  <=  1;
            "HEIGHT_17_30_0": value  <=  1;
            "HEIGHT_17_30_1": value  <=  1;
            "HEIGHT_17_31_0": value  <=  13;
            "HEIGHT_17_31_1": value  <=  13;
            "HEIGHT_17_32_0": value  <=  2;
            "HEIGHT_17_32_1": value  <=  1;
            "HEIGHT_17_33_0": value  <=  6;
            "HEIGHT_17_33_1": value  <=  6;
            "HEIGHT_17_34_0": value  <=  3;
            "HEIGHT_17_34_1": value  <=  1;
            "HEIGHT_17_35_0": value  <=  10;
            "HEIGHT_17_35_1": value  <=  5;
            "HEIGHT_17_36_0": value  <=  5;
            "HEIGHT_17_36_1": value  <=  5;
            "HEIGHT_17_37_0": value  <=  3;
            "HEIGHT_17_37_1": value  <=  3;
            "HEIGHT_17_38_0": value  <=  8;
            "HEIGHT_17_38_1": value  <=  8;
            "HEIGHT_17_39_0": value  <=  13;
            "HEIGHT_17_39_1": value  <=  13;
            "HEIGHT_17_40_0": value  <=  12;
            "HEIGHT_17_40_1": value  <=  6;
            "HEIGHT_17_40_2": value  <=  6;
            "HEIGHT_17_41_0": value  <=  8;
            "HEIGHT_17_41_1": value  <=  8;
            "HEIGHT_17_42_0": value  <=  6;
            "HEIGHT_17_42_1": value  <=  6;
            "HEIGHT_17_43_0": value  <=  8;
            "HEIGHT_17_43_1": value  <=  8;
            "HEIGHT_17_44_0": value  <=  6;
            "HEIGHT_17_44_1": value  <=  3;
            "HEIGHT_17_45_0": value  <=  2;
            "HEIGHT_17_45_1": value  <=  1;
            "HEIGHT_17_45_2": value  <=  1;
            "HEIGHT_17_46_0": value  <=  2;
            "HEIGHT_17_46_1": value  <=  2;
            "HEIGHT_17_47_0": value  <=  2;
            "HEIGHT_17_47_1": value  <=  1;
            "HEIGHT_17_47_2": value  <=  1;
            "HEIGHT_17_48_0": value  <=  2;
            "HEIGHT_17_48_1": value  <=  2;
            "HEIGHT_17_49_0": value  <=  2;
            "HEIGHT_17_49_1": value  <=  1;
            "HEIGHT_17_49_2": value  <=  1;
            "HEIGHT_17_50_0": value  <=  8;
            "HEIGHT_17_50_1": value  <=  8;
            "HEIGHT_17_51_0": value  <=  3;
            "HEIGHT_17_51_1": value  <=  1;
            "HEIGHT_17_52_0": value  <=  3;
            "HEIGHT_17_52_1": value  <=  1;
            "HEIGHT_17_53_0": value  <=  3;
            "HEIGHT_17_53_1": value  <=  3;
            "HEIGHT_17_54_0": value  <=  3;
            "HEIGHT_17_54_1": value  <=  1;
            "HEIGHT_17_55_0": value  <=  3;
            "HEIGHT_17_55_1": value  <=  1;
            "HEIGHT_17_56_0": value  <=  3;
            "HEIGHT_17_56_1": value  <=  1;
            "HEIGHT_17_57_0": value  <=  3;
            "HEIGHT_17_57_1": value  <=  1;
            "HEIGHT_17_58_0": value  <=  2;
            "HEIGHT_17_58_1": value  <=  1;
            "HEIGHT_17_59_0": value  <=  4;
            "HEIGHT_17_59_1": value  <=  2;
            "HEIGHT_17_60_0": value  <=  2;
            "HEIGHT_17_60_1": value  <=  1;
            "HEIGHT_17_61_0": value  <=  2;
            "HEIGHT_17_61_1": value  <=  1;
            "HEIGHT_17_61_2": value  <=  1;
            "HEIGHT_17_62_0": value  <=  2;
            "HEIGHT_17_62_1": value  <=  1;
            "HEIGHT_17_63_0": value  <=  9;
            "HEIGHT_17_63_1": value  <=  3;
            "HEIGHT_17_64_0": value  <=  3;
            "HEIGHT_17_64_1": value  <=  1;
            "HEIGHT_17_65_0": value  <=  4;
            "HEIGHT_17_65_1": value  <=  2;
            "HEIGHT_17_66_0": value  <=  4;
            "HEIGHT_17_66_1": value  <=  2;
            "HEIGHT_17_67_0": value  <=  13;
            "HEIGHT_17_67_1": value  <=  13;
            "HEIGHT_17_68_0": value  <=  12;
            "HEIGHT_17_68_1": value  <=  6;
            "HEIGHT_17_68_2": value  <=  6;
            "HEIGHT_17_69_0": value  <=  6;
            "HEIGHT_17_69_1": value  <=  3;
            "HEIGHT_17_69_2": value  <=  3;
            "HEIGHT_17_70_0": value  <=  6;
            "HEIGHT_17_70_1": value  <=  3;
            "HEIGHT_17_70_2": value  <=  3;
            "HEIGHT_17_71_0": value  <=  2;
            "HEIGHT_17_71_1": value  <=  1;
            "HEIGHT_17_72_0": value  <=  2;
            "HEIGHT_17_72_1": value  <=  1;
            "HEIGHT_17_73_0": value  <=  13;
            "HEIGHT_17_73_1": value  <=  13;
            "HEIGHT_17_74_0": value  <=  13;
            "HEIGHT_17_74_1": value  <=  13;
            "HEIGHT_17_75_0": value  <=  6;
            "HEIGHT_17_75_1": value  <=  2;
            "HEIGHT_17_76_0": value  <=  2;
            "HEIGHT_17_76_1": value  <=  1;
            "HEIGHT_17_76_2": value  <=  1;
            "HEIGHT_17_77_0": value  <=  6;
            "HEIGHT_17_77_1": value  <=  3;
            "HEIGHT_17_77_2": value  <=  3;
            "HEIGHT_17_78_0": value  <=  2;
            "HEIGHT_17_78_1": value  <=  1;
            "HEIGHT_17_78_2": value  <=  1;
            "HEIGHT_17_79_0": value  <=  6;
            "HEIGHT_17_79_1": value  <=  3;
            "HEIGHT_17_79_2": value  <=  3;
            "HEIGHT_17_80_0": value  <=  3;
            "HEIGHT_17_80_1": value  <=  1;
            "HEIGHT_17_81_0": value  <=  10;
            "HEIGHT_17_81_1": value  <=  5;
            "HEIGHT_17_82_0": value  <=  10;
            "HEIGHT_17_82_1": value  <=  5;
            "HEIGHT_17_83_0": value  <=  2;
            "HEIGHT_17_83_1": value  <=  2;
            "HEIGHT_17_84_0": value  <=  2;
            "HEIGHT_17_84_1": value  <=  1;
            "HEIGHT_17_85_0": value  <=  3;
            "HEIGHT_17_85_1": value  <=  1;
            "HEIGHT_17_86_0": value  <=  18;
            "HEIGHT_17_86_1": value  <=  9;
            "HEIGHT_17_86_2": value  <=  9;
            "HEIGHT_17_87_0": value  <=  12;
            "HEIGHT_17_87_1": value  <=  6;
            "HEIGHT_17_88_0": value  <=  6;
            "HEIGHT_17_88_1": value  <=  2;
            "HEIGHT_17_89_0": value  <=  3;
            "HEIGHT_17_89_1": value  <=  1;
            "HEIGHT_17_90_0": value  <=  3;
            "HEIGHT_17_90_1": value  <=  1;
            "HEIGHT_17_91_0": value  <=  2;
            "HEIGHT_17_91_1": value  <=  2;
            "HEIGHT_17_92_0": value  <=  2;
            "HEIGHT_17_92_1": value  <=  2;
            "HEIGHT_17_93_0": value  <=  1;
            "HEIGHT_17_93_1": value  <=  1;
            "HEIGHT_17_94_0": value  <=  3;
            "HEIGHT_17_94_1": value  <=  3;
            "HEIGHT_17_95_0": value  <=  6;
            "HEIGHT_17_95_1": value  <=  3;
            "HEIGHT_17_95_2": value  <=  3;
            "HEIGHT_17_96_0": value  <=  6;
            "HEIGHT_17_96_1": value  <=  3;
            "HEIGHT_17_96_2": value  <=  3;
            "HEIGHT_17_97_0": value  <=  10;
            "HEIGHT_17_97_1": value  <=  5;
            "HEIGHT_17_97_2": value  <=  5;
            "HEIGHT_17_98_0": value  <=  4;
            "HEIGHT_17_98_1": value  <=  4;
            "HEIGHT_17_99_0": value  <=  1;
            "HEIGHT_17_99_1": value  <=  1;
            "HEIGHT_17_100_0": value  <=  2;
            "HEIGHT_17_100_1": value  <=  1;
            "HEIGHT_17_100_2": value  <=  1;
            "HEIGHT_17_101_0": value  <=  6;
            "HEIGHT_17_101_1": value  <=  3;
            "HEIGHT_17_102_0": value  <=  6;
            "HEIGHT_17_102_1": value  <=  3;
            "HEIGHT_17_103_0": value  <=  1;
            "HEIGHT_17_103_1": value  <=  1;
            "HEIGHT_17_104_0": value  <=  3;
            "HEIGHT_17_104_1": value  <=  1;
            "HEIGHT_17_105_0": value  <=  4;
            "HEIGHT_17_105_1": value  <=  2;
            "HEIGHT_17_106_0": value  <=  3;
            "HEIGHT_17_106_1": value  <=  1;
            "HEIGHT_17_107_0": value  <=  2;
            "HEIGHT_17_107_1": value  <=  2;
            "HEIGHT_17_108_0": value  <=  2;
            "HEIGHT_17_108_1": value  <=  1;
            "HEIGHT_17_109_0": value  <=  6;
            "HEIGHT_17_109_1": value  <=  3;
            "HEIGHT_17_110_0": value  <=  2;
            "HEIGHT_17_110_1": value  <=  1;
            "HEIGHT_17_110_2": value  <=  1;
            "HEIGHT_17_111_0": value  <=  4;
            "HEIGHT_17_111_1": value  <=  2;
            "HEIGHT_17_111_2": value  <=  2;
            "HEIGHT_17_112_0": value  <=  2;
            "HEIGHT_17_112_1": value  <=  2;
            "HEIGHT_17_113_0": value  <=  2;
            "HEIGHT_17_113_1": value  <=  1;
            "HEIGHT_17_113_2": value  <=  1;
            "HEIGHT_17_114_0": value  <=  2;
            "HEIGHT_17_114_1": value  <=  1;
            "HEIGHT_17_114_2": value  <=  1;
            "HEIGHT_17_115_0": value  <=  2;
            "HEIGHT_17_115_1": value  <=  1;
            "HEIGHT_17_116_0": value  <=  2;
            "HEIGHT_17_116_1": value  <=  1;
            "HEIGHT_17_117_0": value  <=  8;
            "HEIGHT_17_117_1": value  <=  4;
            "HEIGHT_17_117_2": value  <=  4;
            "HEIGHT_17_118_0": value  <=  3;
            "HEIGHT_17_118_1": value  <=  1;
            "HEIGHT_17_119_0": value  <=  2;
            "HEIGHT_17_119_1": value  <=  2;
            "HEIGHT_17_120_0": value  <=  15;
            "HEIGHT_17_120_1": value  <=  15;
            "HEIGHT_17_121_0": value  <=  14;
            "HEIGHT_17_121_1": value  <=  14;
            "HEIGHT_17_122_0": value  <=  3;
            "HEIGHT_17_122_1": value  <=  1;
            "HEIGHT_17_123_0": value  <=  19;
            "HEIGHT_17_123_1": value  <=  19;
            "HEIGHT_17_124_0": value  <=  2;
            "HEIGHT_17_124_1": value  <=  1;
            "HEIGHT_17_125_0": value  <=  5;
            "HEIGHT_17_125_1": value  <=  5;
            "HEIGHT_17_126_0": value  <=  5;
            "HEIGHT_17_126_1": value  <=  5;
            "HEIGHT_17_127_0": value  <=  2;
            "HEIGHT_17_127_1": value  <=  1;
            "HEIGHT_17_127_2": value  <=  1;
            "HEIGHT_17_128_0": value  <=  6;
            "HEIGHT_17_128_1": value  <=  2;
            "HEIGHT_17_129_0": value  <=  2;
            "HEIGHT_17_129_1": value  <=  1;
            "HEIGHT_17_129_2": value  <=  1;
            "HEIGHT_17_130_0": value  <=  10;
            "HEIGHT_17_130_1": value  <=  5;
            "HEIGHT_17_131_0": value  <=  2;
            "HEIGHT_17_131_1": value  <=  1;
            "HEIGHT_17_131_2": value  <=  1;
            "HEIGHT_17_132_0": value  <=  2;
            "HEIGHT_17_132_1": value  <=  1;
            "HEIGHT_17_133_0": value  <=  2;
            "HEIGHT_17_133_1": value  <=  1;
            "HEIGHT_17_133_2": value  <=  1;
            "HEIGHT_17_134_0": value  <=  2;
            "HEIGHT_17_134_1": value  <=  1;
            "HEIGHT_17_134_2": value  <=  1;
            "HEIGHT_17_135_0": value  <=  3;
            "HEIGHT_17_135_1": value  <=  1;
            "HEIGHT_17_136_0": value  <=  3;
            "HEIGHT_17_136_1": value  <=  1;
            "HEIGHT_17_137_0": value  <=  3;
            "HEIGHT_17_137_1": value  <=  1;
            "HEIGHT_17_138_0": value  <=  3;
            "HEIGHT_17_138_1": value  <=  1;
            "HEIGHT_17_139_0": value  <=  3;
            "HEIGHT_17_139_1": value  <=  1;
            "HEIGHT_17_140_0": value  <=  3;
            "HEIGHT_17_140_1": value  <=  1;
            "HEIGHT_17_141_0": value  <=  3;
            "HEIGHT_17_141_1": value  <=  1;
            "HEIGHT_17_142_0": value  <=  8;
            "HEIGHT_17_142_1": value  <=  4;
            "HEIGHT_17_142_2": value  <=  4;
            "HEIGHT_17_143_0": value  <=  2;
            "HEIGHT_17_143_1": value  <=  1;
            "HEIGHT_17_143_2": value  <=  1;
            "HEIGHT_17_144_0": value  <=  4;
            "HEIGHT_17_144_1": value  <=  4;
            "HEIGHT_17_145_0": value  <=  3;
            "HEIGHT_17_145_1": value  <=  1;
            "HEIGHT_17_146_0": value  <=  6;
            "HEIGHT_17_146_1": value  <=  2;
            "HEIGHT_17_147_0": value  <=  4;
            "HEIGHT_17_147_1": value  <=  4;
            "HEIGHT_17_148_0": value  <=  6;
            "HEIGHT_17_148_1": value  <=  6;
            "HEIGHT_17_149_0": value  <=  2;
            "HEIGHT_17_149_1": value  <=  2;
            "HEIGHT_17_150_0": value  <=  2;
            "HEIGHT_17_150_1": value  <=  2;
            "HEIGHT_17_151_0": value  <=  13;
            "HEIGHT_17_151_1": value  <=  13;
            "HEIGHT_17_152_0": value  <=  13;
            "HEIGHT_17_152_1": value  <=  13;
            "HEIGHT_17_153_0": value  <=  9;
            "HEIGHT_17_153_1": value  <=  3;
            "HEIGHT_17_154_0": value  <=  12;
            "HEIGHT_17_154_1": value  <=  6;
            "HEIGHT_17_155_0": value  <=  2;
            "HEIGHT_17_155_1": value  <=  1;
            "HEIGHT_17_155_2": value  <=  1;
            "HEIGHT_17_156_0": value  <=  2;
            "HEIGHT_17_156_1": value  <=  1;
            "HEIGHT_17_156_2": value  <=  1;
            "HEIGHT_17_157_0": value  <=  2;
            "HEIGHT_17_157_1": value  <=  1;
            "HEIGHT_17_157_2": value  <=  1;
            "HEIGHT_17_158_0": value  <=  2;
            "HEIGHT_17_158_1": value  <=  1;
            "HEIGHT_17_158_2": value  <=  1;
            "HEIGHT_17_159_0": value  <=  2;
            "HEIGHT_17_159_1": value  <=  1;
            "HEIGHT_18_0_0": value  <=  4;
            "HEIGHT_18_0_1": value  <=  2;
            "HEIGHT_18_1_0": value  <=  1;
            "HEIGHT_18_1_1": value  <=  1;
            "HEIGHT_18_2_0": value  <=  12;
            "HEIGHT_18_2_1": value  <=  6;
            "HEIGHT_18_3_0": value  <=  1;
            "HEIGHT_18_3_1": value  <=  1;
            "HEIGHT_18_4_0": value  <=  4;
            "HEIGHT_18_4_1": value  <=  2;
            "HEIGHT_18_4_2": value  <=  2;
            "HEIGHT_18_5_0": value  <=  13;
            "HEIGHT_18_5_1": value  <=  13;
            "HEIGHT_18_6_0": value  <=  13;
            "HEIGHT_18_6_1": value  <=  13;
            "HEIGHT_18_7_0": value  <=  8;
            "HEIGHT_18_7_1": value  <=  4;
            "HEIGHT_18_8_0": value  <=  5;
            "HEIGHT_18_8_1": value  <=  5;
            "HEIGHT_18_9_0": value  <=  1;
            "HEIGHT_18_9_1": value  <=  1;
            "HEIGHT_18_10_0": value  <=  1;
            "HEIGHT_18_10_1": value  <=  1;
            "HEIGHT_18_11_0": value  <=  10;
            "HEIGHT_18_11_1": value  <=  10;
            "HEIGHT_18_12_0": value  <=  3;
            "HEIGHT_18_12_1": value  <=  1;
            "HEIGHT_18_13_0": value  <=  1;
            "HEIGHT_18_13_1": value  <=  1;
            "HEIGHT_18_14_0": value  <=  2;
            "HEIGHT_18_14_1": value  <=  1;
            "HEIGHT_18_15_0": value  <=  2;
            "HEIGHT_18_15_1": value  <=  1;
            "HEIGHT_18_16_0": value  <=  6;
            "HEIGHT_18_16_1": value  <=  3;
            "HEIGHT_18_17_0": value  <=  4;
            "HEIGHT_18_17_1": value  <=  4;
            "HEIGHT_18_18_0": value  <=  4;
            "HEIGHT_18_18_1": value  <=  4;
            "HEIGHT_18_19_0": value  <=  4;
            "HEIGHT_18_19_1": value  <=  4;
            "HEIGHT_18_20_0": value  <=  3;
            "HEIGHT_18_20_1": value  <=  1;
            "HEIGHT_18_21_0": value  <=  4;
            "HEIGHT_18_21_1": value  <=  4;
            "HEIGHT_18_22_0": value  <=  17;
            "HEIGHT_18_22_1": value  <=  17;
            "HEIGHT_18_23_0": value  <=  1;
            "HEIGHT_18_23_1": value  <=  1;
            "HEIGHT_18_24_0": value  <=  4;
            "HEIGHT_18_24_1": value  <=  4;
            "HEIGHT_18_25_0": value  <=  3;
            "HEIGHT_18_25_1": value  <=  1;
            "HEIGHT_18_26_0": value  <=  3;
            "HEIGHT_18_26_1": value  <=  3;
            "HEIGHT_18_27_0": value  <=  10;
            "HEIGHT_18_27_1": value  <=  5;
            "HEIGHT_18_28_0": value  <=  8;
            "HEIGHT_18_28_1": value  <=  4;
            "HEIGHT_18_29_0": value  <=  2;
            "HEIGHT_18_29_1": value  <=  1;
            "HEIGHT_18_30_0": value  <=  2;
            "HEIGHT_18_30_1": value  <=  1;
            "HEIGHT_18_31_0": value  <=  6;
            "HEIGHT_18_31_1": value  <=  3;
            "HEIGHT_18_32_0": value  <=  6;
            "HEIGHT_18_32_1": value  <=  3;
            "HEIGHT_18_33_0": value  <=  3;
            "HEIGHT_18_33_1": value  <=  1;
            "HEIGHT_18_34_0": value  <=  3;
            "HEIGHT_18_34_1": value  <=  1;
            "HEIGHT_18_35_0": value  <=  6;
            "HEIGHT_18_35_1": value  <=  3;
            "HEIGHT_18_35_2": value  <=  3;
            "HEIGHT_18_36_0": value  <=  2;
            "HEIGHT_18_36_1": value  <=  1;
            "HEIGHT_18_37_0": value  <=  2;
            "HEIGHT_18_37_1": value  <=  1;
            "HEIGHT_18_37_2": value  <=  1;
            "HEIGHT_18_38_0": value  <=  8;
            "HEIGHT_18_38_1": value  <=  4;
            "HEIGHT_18_39_0": value  <=  10;
            "HEIGHT_18_39_1": value  <=  5;
            "HEIGHT_18_39_2": value  <=  5;
            "HEIGHT_18_40_0": value  <=  10;
            "HEIGHT_18_40_1": value  <=  5;
            "HEIGHT_18_40_2": value  <=  5;
            "HEIGHT_18_41_0": value  <=  6;
            "HEIGHT_18_41_1": value  <=  2;
            "HEIGHT_18_42_0": value  <=  2;
            "HEIGHT_18_42_1": value  <=  2;
            "HEIGHT_18_43_0": value  <=  6;
            "HEIGHT_18_43_1": value  <=  2;
            "HEIGHT_18_44_0": value  <=  2;
            "HEIGHT_18_44_1": value  <=  1;
            "HEIGHT_18_44_2": value  <=  1;
            "HEIGHT_18_45_0": value  <=  4;
            "HEIGHT_18_45_1": value  <=  4;
            "HEIGHT_18_46_0": value  <=  2;
            "HEIGHT_18_46_1": value  <=  1;
            "HEIGHT_18_47_0": value  <=  4;
            "HEIGHT_18_47_1": value  <=  4;
            "HEIGHT_18_48_0": value  <=  1;
            "HEIGHT_18_48_1": value  <=  1;
            "HEIGHT_18_49_0": value  <=  3;
            "HEIGHT_18_49_1": value  <=  1;
            "HEIGHT_18_50_0": value  <=  2;
            "HEIGHT_18_50_1": value  <=  2;
            "HEIGHT_18_51_0": value  <=  2;
            "HEIGHT_18_51_1": value  <=  1;
            "HEIGHT_18_52_0": value  <=  2;
            "HEIGHT_18_52_1": value  <=  1;
            "HEIGHT_18_53_0": value  <=  3;
            "HEIGHT_18_53_1": value  <=  1;
            "HEIGHT_18_54_0": value  <=  2;
            "HEIGHT_18_54_1": value  <=  1;
            "HEIGHT_18_55_0": value  <=  3;
            "HEIGHT_18_55_1": value  <=  1;
            "HEIGHT_18_56_0": value  <=  3;
            "HEIGHT_18_56_1": value  <=  1;
            "HEIGHT_18_57_0": value  <=  2;
            "HEIGHT_18_57_1": value  <=  2;
            "HEIGHT_18_58_0": value  <=  3;
            "HEIGHT_18_58_1": value  <=  1;
            "HEIGHT_18_59_0": value  <=  3;
            "HEIGHT_18_59_1": value  <=  1;
            "HEIGHT_18_60_0": value  <=  6;
            "HEIGHT_18_60_1": value  <=  2;
            "HEIGHT_18_61_0": value  <=  6;
            "HEIGHT_18_61_1": value  <=  3;
            "HEIGHT_18_61_2": value  <=  3;
            "HEIGHT_18_62_0": value  <=  4;
            "HEIGHT_18_62_1": value  <=  4;
            "HEIGHT_18_63_0": value  <=  2;
            "HEIGHT_18_63_1": value  <=  2;
            "HEIGHT_18_64_0": value  <=  11;
            "HEIGHT_18_64_1": value  <=  11;
            "HEIGHT_18_65_0": value  <=  6;
            "HEIGHT_18_65_1": value  <=  6;
            "HEIGHT_18_66_0": value  <=  1;
            "HEIGHT_18_66_1": value  <=  1;
            "HEIGHT_18_67_0": value  <=  10;
            "HEIGHT_18_67_1": value  <=  5;
            "HEIGHT_18_67_2": value  <=  5;
            "HEIGHT_18_68_0": value  <=  3;
            "HEIGHT_18_68_1": value  <=  1;
            "HEIGHT_18_69_0": value  <=  3;
            "HEIGHT_18_69_1": value  <=  1;
            "HEIGHT_18_70_0": value  <=  10;
            "HEIGHT_18_70_1": value  <=  5;
            "HEIGHT_18_70_2": value  <=  5;
            "HEIGHT_18_71_0": value  <=  6;
            "HEIGHT_18_71_1": value  <=  2;
            "HEIGHT_18_72_0": value  <=  3;
            "HEIGHT_18_72_1": value  <=  1;
            "HEIGHT_18_73_0": value  <=  2;
            "HEIGHT_18_73_1": value  <=  1;
            "HEIGHT_18_74_0": value  <=  6;
            "HEIGHT_18_74_1": value  <=  2;
            "HEIGHT_18_75_0": value  <=  1;
            "HEIGHT_18_75_1": value  <=  1;
            "HEIGHT_18_76_0": value  <=  6;
            "HEIGHT_18_76_1": value  <=  6;
            "HEIGHT_18_77_0": value  <=  14;
            "HEIGHT_18_77_1": value  <=  14;
            "HEIGHT_18_78_0": value  <=  3;
            "HEIGHT_18_78_1": value  <=  3;
            "HEIGHT_18_79_0": value  <=  2;
            "HEIGHT_18_79_1": value  <=  2;
            "HEIGHT_18_80_0": value  <=  2;
            "HEIGHT_18_80_1": value  <=  2;
            "HEIGHT_18_81_0": value  <=  5;
            "HEIGHT_18_81_1": value  <=  5;
            "HEIGHT_18_82_0": value  <=  5;
            "HEIGHT_18_82_1": value  <=  5;
            "HEIGHT_18_83_0": value  <=  10;
            "HEIGHT_18_83_1": value  <=  10;
            "HEIGHT_18_84_0": value  <=  2;
            "HEIGHT_18_84_1": value  <=  1;
            "HEIGHT_18_85_0": value  <=  6;
            "HEIGHT_18_85_1": value  <=  6;
            "HEIGHT_18_86_0": value  <=  10;
            "HEIGHT_18_86_1": value  <=  5;
            "HEIGHT_18_87_0": value  <=  10;
            "HEIGHT_18_87_1": value  <=  10;
            "HEIGHT_18_88_0": value  <=  3;
            "HEIGHT_18_88_1": value  <=  1;
            "HEIGHT_18_89_0": value  <=  7;
            "HEIGHT_18_89_1": value  <=  7;
            "HEIGHT_18_90_0": value  <=  10;
            "HEIGHT_18_90_1": value  <=  10;
            "HEIGHT_18_91_0": value  <=  7;
            "HEIGHT_18_91_1": value  <=  7;
            "HEIGHT_18_92_0": value  <=  2;
            "HEIGHT_18_92_1": value  <=  1;
            "HEIGHT_18_93_0": value  <=  10;
            "HEIGHT_18_93_1": value  <=  10;
            "HEIGHT_18_94_0": value  <=  10;
            "HEIGHT_18_94_1": value  <=  10;
            "HEIGHT_18_95_0": value  <=  4;
            "HEIGHT_18_95_1": value  <=  4;
            "HEIGHT_18_96_0": value  <=  3;
            "HEIGHT_18_96_1": value  <=  3;
            "HEIGHT_18_97_0": value  <=  6;
            "HEIGHT_18_97_1": value  <=  3;
            "HEIGHT_18_97_2": value  <=  3;
            "HEIGHT_18_98_0": value  <=  6;
            "HEIGHT_18_98_1": value  <=  3;
            "HEIGHT_18_98_2": value  <=  3;
            "HEIGHT_18_99_0": value  <=  7;
            "HEIGHT_18_99_1": value  <=  7;
            "HEIGHT_18_100_0": value  <=  7;
            "HEIGHT_18_100_1": value  <=  7;
            "HEIGHT_18_101_0": value  <=  16;
            "HEIGHT_18_101_1": value  <=  16;
            "HEIGHT_18_102_0": value  <=  16;
            "HEIGHT_18_102_1": value  <=  16;
            "HEIGHT_18_103_0": value  <=  8;
            "HEIGHT_18_103_1": value  <=  4;
            "HEIGHT_18_103_2": value  <=  4;
            "HEIGHT_18_104_0": value  <=  3;
            "HEIGHT_18_104_1": value  <=  1;
            "HEIGHT_18_105_0": value  <=  3;
            "HEIGHT_18_105_1": value  <=  3;
            "HEIGHT_18_106_0": value  <=  3;
            "HEIGHT_18_106_1": value  <=  1;
            "HEIGHT_18_107_0": value  <=  4;
            "HEIGHT_18_107_1": value  <=  4;
            "HEIGHT_18_108_0": value  <=  1;
            "HEIGHT_18_108_1": value  <=  1;
            "HEIGHT_18_109_0": value  <=  9;
            "HEIGHT_18_109_1": value  <=  3;
            "HEIGHT_18_110_0": value  <=  4;
            "HEIGHT_18_110_1": value  <=  2;
            "HEIGHT_18_110_2": value  <=  2;
            "HEIGHT_18_111_0": value  <=  2;
            "HEIGHT_18_111_1": value  <=  1;
            "HEIGHT_18_112_0": value  <=  3;
            "HEIGHT_18_112_1": value  <=  1;
            "HEIGHT_18_113_0": value  <=  10;
            "HEIGHT_18_113_1": value  <=  5;
            "HEIGHT_18_113_2": value  <=  5;
            "HEIGHT_18_114_0": value  <=  2;
            "HEIGHT_18_114_1": value  <=  1;
            "HEIGHT_18_115_0": value  <=  1;
            "HEIGHT_18_115_1": value  <=  1;
            "HEIGHT_18_116_0": value  <=  6;
            "HEIGHT_18_116_1": value  <=  2;
            "HEIGHT_18_117_0": value  <=  3;
            "HEIGHT_18_117_1": value  <=  1;
            "HEIGHT_18_118_0": value  <=  2;
            "HEIGHT_18_118_1": value  <=  1;
            "HEIGHT_18_119_0": value  <=  6;
            "HEIGHT_18_119_1": value  <=  2;
            "HEIGHT_18_120_0": value  <=  1;
            "HEIGHT_18_120_1": value  <=  1;
            "HEIGHT_18_121_0": value  <=  1;
            "HEIGHT_18_121_1": value  <=  1;
            "HEIGHT_18_122_0": value  <=  1;
            "HEIGHT_18_122_1": value  <=  1;
            "HEIGHT_18_123_0": value  <=  4;
            "HEIGHT_18_123_1": value  <=  4;
            "HEIGHT_18_124_0": value  <=  3;
            "HEIGHT_18_124_1": value  <=  3;
            "HEIGHT_18_125_0": value  <=  8;
            "HEIGHT_18_125_1": value  <=  4;
            "HEIGHT_18_126_0": value  <=  2;
            "HEIGHT_18_126_1": value  <=  1;
            "HEIGHT_18_127_0": value  <=  6;
            "HEIGHT_18_127_1": value  <=  2;
            "HEIGHT_18_128_0": value  <=  4;
            "HEIGHT_18_128_1": value  <=  4;
            "HEIGHT_18_129_0": value  <=  6;
            "HEIGHT_18_129_1": value  <=  2;
            "HEIGHT_18_130_0": value  <=  1;
            "HEIGHT_18_130_1": value  <=  1;
            "HEIGHT_18_131_0": value  <=  4;
            "HEIGHT_18_131_1": value  <=  4;
            "HEIGHT_18_132_0": value  <=  4;
            "HEIGHT_18_132_1": value  <=  2;
            "HEIGHT_18_133_0": value  <=  4;
            "HEIGHT_18_133_1": value  <=  4;
            "HEIGHT_18_134_0": value  <=  4;
            "HEIGHT_18_134_1": value  <=  4;
            "HEIGHT_18_135_0": value  <=  3;
            "HEIGHT_18_135_1": value  <=  1;
            "HEIGHT_18_136_0": value  <=  6;
            "HEIGHT_18_136_1": value  <=  3;
            "HEIGHT_18_137_0": value  <=  12;
            "HEIGHT_18_137_1": value  <=  4;
            "HEIGHT_18_138_0": value  <=  3;
            "HEIGHT_18_138_1": value  <=  1;
            "HEIGHT_18_139_0": value  <=  2;
            "HEIGHT_18_139_1": value  <=  1;
            "HEIGHT_18_139_2": value  <=  1;
            "HEIGHT_18_140_0": value  <=  2;
            "HEIGHT_18_140_1": value  <=  1;
            "HEIGHT_18_141_0": value  <=  15;
            "HEIGHT_18_141_1": value  <=  15;
            "HEIGHT_18_142_0": value  <=  2;
            "HEIGHT_18_142_1": value  <=  1;
            "HEIGHT_18_143_0": value  <=  3;
            "HEIGHT_18_143_1": value  <=  3;
            "HEIGHT_18_144_0": value  <=  15;
            "HEIGHT_18_144_1": value  <=  15;
            "HEIGHT_18_145_0": value  <=  8;
            "HEIGHT_18_145_1": value  <=  4;
            "HEIGHT_18_145_2": value  <=  4;
            "HEIGHT_18_146_0": value  <=  16;
            "HEIGHT_18_146_1": value  <=  8;
            "HEIGHT_18_146_2": value  <=  8;
            "HEIGHT_18_147_0": value  <=  12;
            "HEIGHT_18_147_1": value  <=  6;
            "HEIGHT_18_148_0": value  <=  12;
            "HEIGHT_18_148_1": value  <=  6;
            "HEIGHT_18_148_2": value  <=  6;
            "HEIGHT_18_149_0": value  <=  3;
            "HEIGHT_18_149_1": value  <=  1;
            "HEIGHT_18_150_0": value  <=  3;
            "HEIGHT_18_150_1": value  <=  1;
            "HEIGHT_18_151_0": value  <=  10;
            "HEIGHT_18_151_1": value  <=  5;
            "HEIGHT_18_151_2": value  <=  5;
            "HEIGHT_18_152_0": value  <=  3;
            "HEIGHT_18_152_1": value  <=  1;
            "HEIGHT_18_153_0": value  <=  2;
            "HEIGHT_18_153_1": value  <=  1;
            "HEIGHT_18_153_2": value  <=  1;
            "HEIGHT_18_154_0": value  <=  2;
            "HEIGHT_18_154_1": value  <=  1;
            "HEIGHT_18_154_2": value  <=  1;
            "HEIGHT_18_155_0": value  <=  6;
            "HEIGHT_18_155_1": value  <=  3;
            "HEIGHT_18_155_2": value  <=  3;
            "HEIGHT_18_156_0": value  <=  6;
            "HEIGHT_18_156_1": value  <=  3;
            "HEIGHT_18_156_2": value  <=  3;
            "HEIGHT_18_157_0": value  <=  6;
            "HEIGHT_18_157_1": value  <=  3;
            "HEIGHT_18_158_0": value  <=  10;
            "HEIGHT_18_158_1": value  <=  5;
            "HEIGHT_18_158_2": value  <=  5;
            "HEIGHT_18_159_0": value  <=  2;
            "HEIGHT_18_159_1": value  <=  1;
            "HEIGHT_18_159_2": value  <=  1;
            "HEIGHT_18_160_0": value  <=  8;
            "HEIGHT_18_160_1": value  <=  8;
            "HEIGHT_18_161_0": value  <=  10;
            "HEIGHT_18_161_1": value  <=  5;
            "HEIGHT_18_161_2": value  <=  5;
            "HEIGHT_18_162_0": value  <=  1;
            "HEIGHT_18_162_1": value  <=  1;
            "HEIGHT_18_163_0": value  <=  12;
            "HEIGHT_18_163_1": value  <=  4;
            "HEIGHT_18_164_0": value  <=  9;
            "HEIGHT_18_164_1": value  <=  9;
            "HEIGHT_18_165_0": value  <=  10;
            "HEIGHT_18_165_1": value  <=  5;
            "HEIGHT_18_165_2": value  <=  5;
            "HEIGHT_18_166_0": value  <=  10;
            "HEIGHT_18_166_1": value  <=  5;
            "HEIGHT_18_166_2": value  <=  5;
            "HEIGHT_18_167_0": value  <=  2;
            "HEIGHT_18_167_1": value  <=  1;
            "HEIGHT_18_167_2": value  <=  1;
            "HEIGHT_18_168_0": value  <=  3;
            "HEIGHT_18_168_1": value  <=  1;
            "HEIGHT_18_169_0": value  <=  2;
            "HEIGHT_18_169_1": value  <=  1;
            "HEIGHT_18_169_2": value  <=  1;
            "HEIGHT_18_170_0": value  <=  2;
            "HEIGHT_18_170_1": value  <=  2;
            "HEIGHT_18_171_0": value  <=  2;
            "HEIGHT_18_171_1": value  <=  1;
            "HEIGHT_18_171_2": value  <=  1;
            "HEIGHT_18_172_0": value  <=  2;
            "HEIGHT_18_172_1": value  <=  1;
            "HEIGHT_18_172_2": value  <=  1;
            "HEIGHT_18_173_0": value  <=  12;
            "HEIGHT_18_173_1": value  <=  6;
            "HEIGHT_18_173_2": value  <=  6;
            "HEIGHT_18_174_0": value  <=  10;
            "HEIGHT_18_174_1": value  <=  10;
            "HEIGHT_18_175_0": value  <=  8;
            "HEIGHT_18_175_1": value  <=  4;
            "HEIGHT_18_176_0": value  <=  4;
            "HEIGHT_18_176_1": value  <=  2;
            "HEIGHT_19_0_0": value  <=  2;
            "HEIGHT_19_0_1": value  <=  2;
            "HEIGHT_19_1_0": value  <=  3;
            "HEIGHT_19_1_1": value  <=  1;
            "HEIGHT_19_2_0": value  <=  4;
            "HEIGHT_19_2_1": value  <=  2;
            "HEIGHT_19_2_2": value  <=  2;
            "HEIGHT_19_3_0": value  <=  9;
            "HEIGHT_19_3_1": value  <=  3;
            "HEIGHT_19_4_0": value  <=  4;
            "HEIGHT_19_4_1": value  <=  2;
            "HEIGHT_19_5_0": value  <=  7;
            "HEIGHT_19_5_1": value  <=  7;
            "HEIGHT_19_6_0": value  <=  10;
            "HEIGHT_19_6_1": value  <=  5;
            "HEIGHT_19_6_2": value  <=  5;
            "HEIGHT_19_7_0": value  <=  2;
            "HEIGHT_19_7_1": value  <=  1;
            "HEIGHT_19_8_0": value  <=  15;
            "HEIGHT_19_8_1": value  <=  5;
            "HEIGHT_19_9_0": value  <=  2;
            "HEIGHT_19_9_1": value  <=  1;
            "HEIGHT_19_10_0": value  <=  2;
            "HEIGHT_19_10_1": value  <=  2;
            "HEIGHT_19_11_0": value  <=  15;
            "HEIGHT_19_11_1": value  <=  5;
            "HEIGHT_19_12_0": value  <=  6;
            "HEIGHT_19_12_1": value  <=  3;
            "HEIGHT_19_13_0": value  <=  2;
            "HEIGHT_19_13_1": value  <=  2;
            "HEIGHT_19_14_0": value  <=  1;
            "HEIGHT_19_14_1": value  <=  1;
            "HEIGHT_19_15_0": value  <=  3;
            "HEIGHT_19_15_1": value  <=  1;
            "HEIGHT_19_16_0": value  <=  2;
            "HEIGHT_19_16_1": value  <=  1;
            "HEIGHT_19_17_0": value  <=  3;
            "HEIGHT_19_17_1": value  <=  1;
            "HEIGHT_19_18_0": value  <=  1;
            "HEIGHT_19_18_1": value  <=  1;
            "HEIGHT_19_19_0": value  <=  14;
            "HEIGHT_19_19_1": value  <=  7;
            "HEIGHT_19_20_0": value  <=  10;
            "HEIGHT_19_20_1": value  <=  5;
            "HEIGHT_19_20_2": value  <=  5;
            "HEIGHT_19_21_0": value  <=  2;
            "HEIGHT_19_21_1": value  <=  2;
            "HEIGHT_19_22_0": value  <=  2;
            "HEIGHT_19_22_1": value  <=  2;
            "HEIGHT_19_23_0": value  <=  3;
            "HEIGHT_19_23_1": value  <=  1;
            "HEIGHT_19_24_0": value  <=  16;
            "HEIGHT_19_24_1": value  <=  8;
            "HEIGHT_19_25_0": value  <=  3;
            "HEIGHT_19_25_1": value  <=  1;
            "HEIGHT_19_26_0": value  <=  6;
            "HEIGHT_19_26_1": value  <=  2;
            "HEIGHT_19_27_0": value  <=  9;
            "HEIGHT_19_27_1": value  <=  3;
            "HEIGHT_19_28_0": value  <=  3;
            "HEIGHT_19_28_1": value  <=  1;
            "HEIGHT_19_29_0": value  <=  2;
            "HEIGHT_19_29_1": value  <=  2;
            "HEIGHT_19_30_0": value  <=  3;
            "HEIGHT_19_30_1": value  <=  1;
            "HEIGHT_19_31_0": value  <=  6;
            "HEIGHT_19_31_1": value  <=  2;
            "HEIGHT_19_32_0": value  <=  6;
            "HEIGHT_19_32_1": value  <=  3;
            "HEIGHT_19_33_0": value  <=  2;
            "HEIGHT_19_33_1": value  <=  1;
            "HEIGHT_19_34_0": value  <=  2;
            "HEIGHT_19_34_1": value  <=  1;
            "HEIGHT_19_35_0": value  <=  2;
            "HEIGHT_19_35_1": value  <=  1;
            "HEIGHT_19_36_0": value  <=  6;
            "HEIGHT_19_36_1": value  <=  2;
            "HEIGHT_19_37_0": value  <=  3;
            "HEIGHT_19_37_1": value  <=  1;
            "HEIGHT_19_38_0": value  <=  6;
            "HEIGHT_19_38_1": value  <=  2;
            "HEIGHT_19_39_0": value  <=  3;
            "HEIGHT_19_39_1": value  <=  1;
            "HEIGHT_19_40_0": value  <=  3;
            "HEIGHT_19_40_1": value  <=  1;
            "HEIGHT_19_41_0": value  <=  3;
            "HEIGHT_19_41_1": value  <=  1;
            "HEIGHT_19_42_0": value  <=  12;
            "HEIGHT_19_42_1": value  <=  6;
            "HEIGHT_19_43_0": value  <=  3;
            "HEIGHT_19_43_1": value  <=  1;
            "HEIGHT_19_44_0": value  <=  2;
            "HEIGHT_19_44_1": value  <=  2;
            "HEIGHT_19_45_0": value  <=  3;
            "HEIGHT_19_45_1": value  <=  1;
            "HEIGHT_19_46_0": value  <=  3;
            "HEIGHT_19_46_1": value  <=  1;
            "HEIGHT_19_47_0": value  <=  2;
            "HEIGHT_19_47_1": value  <=  2;
            "HEIGHT_19_48_0": value  <=  3;
            "HEIGHT_19_48_1": value  <=  1;
            "HEIGHT_19_49_0": value  <=  6;
            "HEIGHT_19_49_1": value  <=  6;
            "HEIGHT_19_50_0": value  <=  7;
            "HEIGHT_19_50_1": value  <=  7;
            "HEIGHT_19_51_0": value  <=  3;
            "HEIGHT_19_51_1": value  <=  3;
            "HEIGHT_19_52_0": value  <=  3;
            "HEIGHT_19_52_1": value  <=  3;
            "HEIGHT_19_53_0": value  <=  3;
            "HEIGHT_19_53_1": value  <=  1;
            "HEIGHT_19_54_0": value  <=  1;
            "HEIGHT_19_54_1": value  <=  1;
            "HEIGHT_19_55_0": value  <=  2;
            "HEIGHT_19_55_1": value  <=  2;
            "HEIGHT_19_56_0": value  <=  2;
            "HEIGHT_19_56_1": value  <=  2;
            "HEIGHT_19_57_0": value  <=  2;
            "HEIGHT_19_57_1": value  <=  2;
            "HEIGHT_19_58_0": value  <=  2;
            "HEIGHT_19_58_1": value  <=  2;
            "HEIGHT_19_59_0": value  <=  4;
            "HEIGHT_19_59_1": value  <=  2;
            "HEIGHT_19_60_0": value  <=  2;
            "HEIGHT_19_60_1": value  <=  2;
            "HEIGHT_19_61_0": value  <=  3;
            "HEIGHT_19_61_1": value  <=  1;
            "HEIGHT_19_62_0": value  <=  12;
            "HEIGHT_19_62_1": value  <=  6;
            "HEIGHT_19_62_2": value  <=  6;
            "HEIGHT_19_63_0": value  <=  8;
            "HEIGHT_19_63_1": value  <=  4;
            "HEIGHT_19_63_2": value  <=  4;
            "HEIGHT_19_64_0": value  <=  4;
            "HEIGHT_19_64_1": value  <=  4;
            "HEIGHT_19_65_0": value  <=  1;
            "HEIGHT_19_65_1": value  <=  1;
            "HEIGHT_19_66_0": value  <=  2;
            "HEIGHT_19_66_1": value  <=  1;
            "HEIGHT_19_67_0": value  <=  3;
            "HEIGHT_19_67_1": value  <=  1;
            "HEIGHT_19_68_0": value  <=  3;
            "HEIGHT_19_68_1": value  <=  1;
            "HEIGHT_19_69_0": value  <=  3;
            "HEIGHT_19_69_1": value  <=  1;
            "HEIGHT_19_70_0": value  <=  4;
            "HEIGHT_19_70_1": value  <=  2;
            "HEIGHT_19_70_2": value  <=  2;
            "HEIGHT_19_71_0": value  <=  2;
            "HEIGHT_19_71_1": value  <=  1;
            "HEIGHT_19_71_2": value  <=  1;
            "HEIGHT_19_72_0": value  <=  2;
            "HEIGHT_19_72_1": value  <=  2;
            "HEIGHT_19_73_0": value  <=  2;
            "HEIGHT_19_73_1": value  <=  1;
            "HEIGHT_19_73_2": value  <=  1;
            "HEIGHT_19_74_0": value  <=  3;
            "HEIGHT_19_74_1": value  <=  1;
            "HEIGHT_19_75_0": value  <=  2;
            "HEIGHT_19_75_1": value  <=  1;
            "HEIGHT_19_75_2": value  <=  1;
            "HEIGHT_19_76_0": value  <=  2;
            "HEIGHT_19_76_1": value  <=  1;
            "HEIGHT_19_76_2": value  <=  1;
            "HEIGHT_19_77_0": value  <=  4;
            "HEIGHT_19_77_1": value  <=  4;
            "HEIGHT_19_78_0": value  <=  4;
            "HEIGHT_19_78_1": value  <=  4;
            "HEIGHT_19_79_0": value  <=  1;
            "HEIGHT_19_79_1": value  <=  1;
            "HEIGHT_19_80_0": value  <=  1;
            "HEIGHT_19_80_1": value  <=  1;
            "HEIGHT_19_81_0": value  <=  2;
            "HEIGHT_19_81_1": value  <=  1;
            "HEIGHT_19_81_2": value  <=  1;
            "HEIGHT_19_82_0": value  <=  1;
            "HEIGHT_19_82_1": value  <=  1;
            "HEIGHT_19_83_0": value  <=  8;
            "HEIGHT_19_83_1": value  <=  4;
            "HEIGHT_19_83_2": value  <=  4;
            "HEIGHT_19_84_0": value  <=  2;
            "HEIGHT_19_84_1": value  <=  1;
            "HEIGHT_19_85_0": value  <=  2;
            "HEIGHT_19_85_1": value  <=  1;
            "HEIGHT_19_86_0": value  <=  12;
            "HEIGHT_19_86_1": value  <=  6;
            "HEIGHT_19_86_2": value  <=  6;
            "HEIGHT_19_87_0": value  <=  3;
            "HEIGHT_19_87_1": value  <=  1;
            "HEIGHT_19_88_0": value  <=  2;
            "HEIGHT_19_88_1": value  <=  2;
            "HEIGHT_19_89_0": value  <=  1;
            "HEIGHT_19_89_1": value  <=  1;
            "HEIGHT_19_90_0": value  <=  1;
            "HEIGHT_19_90_1": value  <=  1;
            "HEIGHT_19_91_0": value  <=  2;
            "HEIGHT_19_91_1": value  <=  1;
            "HEIGHT_19_91_2": value  <=  1;
            "HEIGHT_19_92_0": value  <=  3;
            "HEIGHT_19_92_1": value  <=  1;
            "HEIGHT_19_93_0": value  <=  3;
            "HEIGHT_19_93_1": value  <=  3;
            "HEIGHT_19_94_0": value  <=  14;
            "HEIGHT_19_94_1": value  <=  14;
            "HEIGHT_19_95_0": value  <=  3;
            "HEIGHT_19_95_1": value  <=  3;
            "HEIGHT_19_96_0": value  <=  3;
            "HEIGHT_19_96_1": value  <=  3;
            "HEIGHT_19_97_0": value  <=  6;
            "HEIGHT_19_97_1": value  <=  3;
            "HEIGHT_19_98_0": value  <=  8;
            "HEIGHT_19_98_1": value  <=  4;
            "HEIGHT_19_99_0": value  <=  3;
            "HEIGHT_19_99_1": value  <=  1;
            "HEIGHT_19_100_0": value  <=  12;
            "HEIGHT_19_100_1": value  <=  4;
            "HEIGHT_19_101_0": value  <=  3;
            "HEIGHT_19_101_1": value  <=  1;
            "HEIGHT_19_102_0": value  <=  8;
            "HEIGHT_19_102_1": value  <=  8;
            "HEIGHT_19_103_0": value  <=  2;
            "HEIGHT_19_103_1": value  <=  1;
            "HEIGHT_19_103_2": value  <=  1;
            "HEIGHT_19_104_0": value  <=  14;
            "HEIGHT_19_104_1": value  <=  7;
            "HEIGHT_19_105_0": value  <=  2;
            "HEIGHT_19_105_1": value  <=  1;
            "HEIGHT_19_105_2": value  <=  1;
            "HEIGHT_19_106_0": value  <=  2;
            "HEIGHT_19_106_1": value  <=  1;
            "HEIGHT_19_106_2": value  <=  1;
            "HEIGHT_19_107_0": value  <=  3;
            "HEIGHT_19_107_1": value  <=  1;
            "HEIGHT_19_108_0": value  <=  3;
            "HEIGHT_19_108_1": value  <=  1;
            "HEIGHT_19_109_0": value  <=  3;
            "HEIGHT_19_109_1": value  <=  1;
            "HEIGHT_19_110_0": value  <=  3;
            "HEIGHT_19_110_1": value  <=  1;
            "HEIGHT_19_111_0": value  <=  2;
            "HEIGHT_19_111_1": value  <=  1;
            "HEIGHT_19_112_0": value  <=  2;
            "HEIGHT_19_112_1": value  <=  1;
            "HEIGHT_19_112_2": value  <=  1;
            "HEIGHT_19_113_0": value  <=  3;
            "HEIGHT_19_113_1": value  <=  1;
            "HEIGHT_19_114_0": value  <=  2;
            "HEIGHT_19_114_1": value  <=  1;
            "HEIGHT_19_115_0": value  <=  9;
            "HEIGHT_19_115_1": value  <=  3;
            "HEIGHT_19_116_0": value  <=  3;
            "HEIGHT_19_116_1": value  <=  3;
            "HEIGHT_19_117_0": value  <=  3;
            "HEIGHT_19_117_1": value  <=  1;
            "HEIGHT_19_118_0": value  <=  9;
            "HEIGHT_19_118_1": value  <=  3;
            "HEIGHT_19_119_0": value  <=  6;
            "HEIGHT_19_119_1": value  <=  6;
            "HEIGHT_19_120_0": value  <=  6;
            "HEIGHT_19_120_1": value  <=  6;
            "HEIGHT_19_121_0": value  <=  2;
            "HEIGHT_19_121_1": value  <=  1;
            "HEIGHT_19_122_0": value  <=  3;
            "HEIGHT_19_122_1": value  <=  3;
            "HEIGHT_19_123_0": value  <=  3;
            "HEIGHT_19_123_1": value  <=  1;
            "HEIGHT_19_124_0": value  <=  3;
            "HEIGHT_19_124_1": value  <=  1;
            "HEIGHT_19_125_0": value  <=  8;
            "HEIGHT_19_125_1": value  <=  4;
            "HEIGHT_19_125_2": value  <=  4;
            "HEIGHT_19_126_0": value  <=  8;
            "HEIGHT_19_126_1": value  <=  4;
            "HEIGHT_19_126_2": value  <=  4;
            "HEIGHT_19_127_0": value  <=  6;
            "HEIGHT_19_127_1": value  <=  3;
            "HEIGHT_19_128_0": value  <=  20;
            "HEIGHT_19_128_1": value  <=  20;
            "HEIGHT_19_129_0": value  <=  2;
            "HEIGHT_19_129_1": value  <=  2;
            "HEIGHT_19_130_0": value  <=  2;
            "HEIGHT_19_130_1": value  <=  2;
            "HEIGHT_19_131_0": value  <=  1;
            "HEIGHT_19_131_1": value  <=  1;
            "HEIGHT_19_132_0": value  <=  3;
            "HEIGHT_19_132_1": value  <=  3;
            "HEIGHT_19_133_0": value  <=  5;
            "HEIGHT_19_133_1": value  <=  5;
            "HEIGHT_19_134_0": value  <=  2;
            "HEIGHT_19_134_1": value  <=  2;
            "HEIGHT_19_135_0": value  <=  15;
            "HEIGHT_19_135_1": value  <=  15;
            "HEIGHT_19_136_0": value  <=  1;
            "HEIGHT_19_136_1": value  <=  1;
            "HEIGHT_19_137_0": value  <=  4;
            "HEIGHT_19_137_1": value  <=  4;
            "HEIGHT_19_138_0": value  <=  1;
            "HEIGHT_19_138_1": value  <=  1;
            "HEIGHT_19_139_0": value  <=  2;
            "HEIGHT_19_139_1": value  <=  1;
            "HEIGHT_19_140_0": value  <=  6;
            "HEIGHT_19_140_1": value  <=  3;
            "HEIGHT_19_141_0": value  <=  2;
            "HEIGHT_19_141_1": value  <=  1;
            "HEIGHT_19_142_0": value  <=  3;
            "HEIGHT_19_142_1": value  <=  1;
            "HEIGHT_19_143_0": value  <=  10;
            "HEIGHT_19_143_1": value  <=  5;
            "HEIGHT_19_143_2": value  <=  5;
            "HEIGHT_19_144_0": value  <=  2;
            "HEIGHT_19_144_1": value  <=  1;
            "HEIGHT_19_145_0": value  <=  2;
            "HEIGHT_19_145_1": value  <=  1;
            "HEIGHT_19_145_2": value  <=  1;
            "HEIGHT_19_146_0": value  <=  3;
            "HEIGHT_19_146_1": value  <=  1;
            "HEIGHT_19_147_0": value  <=  2;
            "HEIGHT_19_147_1": value  <=  1;
            "HEIGHT_19_148_0": value  <=  2;
            "HEIGHT_19_148_1": value  <=  1;
            "HEIGHT_19_149_0": value  <=  9;
            "HEIGHT_19_149_1": value  <=  3;
            "HEIGHT_19_150_0": value  <=  7;
            "HEIGHT_19_150_1": value  <=  7;
            "HEIGHT_19_151_0": value  <=  5;
            "HEIGHT_19_151_1": value  <=  5;
            "HEIGHT_19_152_0": value  <=  2;
            "HEIGHT_19_152_1": value  <=  1;
            "HEIGHT_19_152_2": value  <=  1;
            "HEIGHT_19_153_0": value  <=  2;
            "HEIGHT_19_153_1": value  <=  1;
            "HEIGHT_19_154_0": value  <=  2;
            "HEIGHT_19_154_1": value  <=  1;
            "HEIGHT_19_155_0": value  <=  8;
            "HEIGHT_19_155_1": value  <=  4;
            "HEIGHT_19_155_2": value  <=  4;
            "HEIGHT_19_156_0": value  <=  6;
            "HEIGHT_19_156_1": value  <=  6;
            "HEIGHT_19_157_0": value  <=  17;
            "HEIGHT_19_157_1": value  <=  17;
            "HEIGHT_19_158_0": value  <=  1;
            "HEIGHT_19_158_1": value  <=  1;
            "HEIGHT_19_159_0": value  <=  5;
            "HEIGHT_19_159_1": value  <=  5;
            "HEIGHT_19_160_0": value  <=  5;
            "HEIGHT_19_160_1": value  <=  5;
            "HEIGHT_19_161_0": value  <=  4;
            "HEIGHT_19_161_1": value  <=  2;
            "HEIGHT_19_161_2": value  <=  2;
            "HEIGHT_19_162_0": value  <=  2;
            "HEIGHT_19_162_1": value  <=  1;
            "HEIGHT_19_162_2": value  <=  1;
            "HEIGHT_19_163_0": value  <=  3;
            "HEIGHT_19_163_1": value  <=  1;
            "HEIGHT_19_164_0": value  <=  2;
            "HEIGHT_19_164_1": value  <=  1;
            "HEIGHT_19_164_2": value  <=  1;
            "HEIGHT_19_165_0": value  <=  8;
            "HEIGHT_19_165_1": value  <=  4;
            "HEIGHT_19_165_2": value  <=  4;
            "HEIGHT_19_166_0": value  <=  6;
            "HEIGHT_19_166_1": value  <=  3;
            "HEIGHT_19_167_0": value  <=  2;
            "HEIGHT_19_167_1": value  <=  1;
            "HEIGHT_19_168_0": value  <=  2;
            "HEIGHT_19_168_1": value  <=  1;
            "HEIGHT_19_168_2": value  <=  1;
            "HEIGHT_19_169_0": value  <=  4;
            "HEIGHT_19_169_1": value  <=  2;
            "HEIGHT_19_169_2": value  <=  2;
            "HEIGHT_19_170_0": value  <=  2;
            "HEIGHT_19_170_1": value  <=  1;
            "HEIGHT_19_171_0": value  <=  3;
            "HEIGHT_19_171_1": value  <=  3;
            "HEIGHT_19_172_0": value  <=  2;
            "HEIGHT_19_172_1": value  <=  1;
            "HEIGHT_19_173_0": value  <=  12;
            "HEIGHT_19_173_1": value  <=  6;
            "HEIGHT_19_173_2": value  <=  6;
            "HEIGHT_19_174_0": value  <=  12;
            "HEIGHT_19_174_1": value  <=  6;
            "HEIGHT_19_174_2": value  <=  6;
            "HEIGHT_19_175_0": value  <=  10;
            "HEIGHT_19_175_1": value  <=  10;
            "HEIGHT_19_176_0": value  <=  4;
            "HEIGHT_19_176_1": value  <=  2;
            "HEIGHT_19_176_2": value  <=  2;
            "HEIGHT_19_177_0": value  <=  4;
            "HEIGHT_19_177_1": value  <=  2;
            "HEIGHT_19_177_2": value  <=  2;
            "HEIGHT_19_178_0": value  <=  6;
            "HEIGHT_19_178_1": value  <=  6;
            "HEIGHT_19_179_0": value  <=  10;
            "HEIGHT_19_179_1": value  <=  10;
            "HEIGHT_19_180_0": value  <=  9;
            "HEIGHT_19_180_1": value  <=  9;
            "HEIGHT_19_181_0": value  <=  1;
            "HEIGHT_19_181_1": value  <=  1;
            "HEIGHT_20_0_0": value  <=  9;
            "HEIGHT_20_0_1": value  <=  9;
            "HEIGHT_20_1_0": value  <=  4;
            "HEIGHT_20_1_1": value  <=  4;
            "HEIGHT_20_2_0": value  <=  4;
            "HEIGHT_20_2_1": value  <=  2;
            "HEIGHT_20_3_0": value  <=  8;
            "HEIGHT_20_3_1": value  <=  4;
            "HEIGHT_20_4_0": value  <=  12;
            "HEIGHT_20_4_1": value  <=  6;
            "HEIGHT_20_5_0": value  <=  6;
            "HEIGHT_20_5_1": value  <=  3;
            "HEIGHT_20_6_0": value  <=  6;
            "HEIGHT_20_6_1": value  <=  3;
            "HEIGHT_20_7_0": value  <=  4;
            "HEIGHT_20_7_1": value  <=  2;
            "HEIGHT_20_7_2": value  <=  2;
            "HEIGHT_20_8_0": value  <=  2;
            "HEIGHT_20_8_1": value  <=  2;
            "HEIGHT_20_9_0": value  <=  2;
            "HEIGHT_20_9_1": value  <=  1;
            "HEIGHT_20_10_0": value  <=  6;
            "HEIGHT_20_10_1": value  <=  2;
            "HEIGHT_20_11_0": value  <=  2;
            "HEIGHT_20_11_1": value  <=  1;
            "HEIGHT_20_12_0": value  <=  3;
            "HEIGHT_20_12_1": value  <=  1;
            "HEIGHT_20_13_0": value  <=  2;
            "HEIGHT_20_13_1": value  <=  1;
            "HEIGHT_20_14_0": value  <=  2;
            "HEIGHT_20_14_1": value  <=  1;
            "HEIGHT_20_15_0": value  <=  7;
            "HEIGHT_20_15_1": value  <=  7;
            "HEIGHT_20_16_0": value  <=  6;
            "HEIGHT_20_16_1": value  <=  2;
            "HEIGHT_20_17_0": value  <=  3;
            "HEIGHT_20_17_1": value  <=  1;
            "HEIGHT_20_18_0": value  <=  2;
            "HEIGHT_20_18_1": value  <=  2;
            "HEIGHT_20_19_0": value  <=  3;
            "HEIGHT_20_19_1": value  <=  1;
            "HEIGHT_20_20_0": value  <=  3;
            "HEIGHT_20_20_1": value  <=  1;
            "HEIGHT_20_21_0": value  <=  2;
            "HEIGHT_20_21_1": value  <=  1;
            "HEIGHT_20_22_0": value  <=  3;
            "HEIGHT_20_22_1": value  <=  3;
            "HEIGHT_20_23_0": value  <=  7;
            "HEIGHT_20_23_1": value  <=  7;
            "HEIGHT_20_24_0": value  <=  1;
            "HEIGHT_20_24_1": value  <=  1;
            "HEIGHT_20_25_0": value  <=  3;
            "HEIGHT_20_25_1": value  <=  1;
            "HEIGHT_20_26_0": value  <=  4;
            "HEIGHT_20_26_1": value  <=  4;
            "HEIGHT_20_27_0": value  <=  6;
            "HEIGHT_20_27_1": value  <=  2;
            "HEIGHT_20_28_0": value  <=  6;
            "HEIGHT_20_28_1": value  <=  2;
            "HEIGHT_20_29_0": value  <=  6;
            "HEIGHT_20_29_1": value  <=  3;
            "HEIGHT_20_29_2": value  <=  3;
            "HEIGHT_20_30_0": value  <=  3;
            "HEIGHT_20_30_1": value  <=  1;
            "HEIGHT_20_31_0": value  <=  6;
            "HEIGHT_20_31_1": value  <=  3;
            "HEIGHT_20_31_2": value  <=  3;
            "HEIGHT_20_32_0": value  <=  3;
            "HEIGHT_20_32_1": value  <=  1;
            "HEIGHT_20_33_0": value  <=  3;
            "HEIGHT_20_33_1": value  <=  1;
            "HEIGHT_20_34_0": value  <=  3;
            "HEIGHT_20_34_1": value  <=  1;
            "HEIGHT_20_35_0": value  <=  3;
            "HEIGHT_20_35_1": value  <=  1;
            "HEIGHT_20_36_0": value  <=  2;
            "HEIGHT_20_36_1": value  <=  1;
            "HEIGHT_20_37_0": value  <=  3;
            "HEIGHT_20_37_1": value  <=  1;
            "HEIGHT_20_38_0": value  <=  4;
            "HEIGHT_20_38_1": value  <=  2;
            "HEIGHT_20_39_0": value  <=  3;
            "HEIGHT_20_39_1": value  <=  3;
            "HEIGHT_20_40_0": value  <=  3;
            "HEIGHT_20_40_1": value  <=  3;
            "HEIGHT_20_41_0": value  <=  6;
            "HEIGHT_20_41_1": value  <=  6;
            "HEIGHT_20_42_0": value  <=  7;
            "HEIGHT_20_42_1": value  <=  7;
            "HEIGHT_20_43_0": value  <=  6;
            "HEIGHT_20_43_1": value  <=  6;
            "HEIGHT_20_44_0": value  <=  3;
            "HEIGHT_20_44_1": value  <=  1;
            "HEIGHT_20_45_0": value  <=  6;
            "HEIGHT_20_45_1": value  <=  6;
            "HEIGHT_20_46_0": value  <=  6;
            "HEIGHT_20_46_1": value  <=  6;
            "HEIGHT_20_47_0": value  <=  1;
            "HEIGHT_20_47_1": value  <=  1;
            "HEIGHT_20_48_0": value  <=  7;
            "HEIGHT_20_48_1": value  <=  7;
            "HEIGHT_20_49_0": value  <=  2;
            "HEIGHT_20_49_1": value  <=  1;
            "HEIGHT_20_50_0": value  <=  2;
            "HEIGHT_20_50_1": value  <=  1;
            "HEIGHT_20_51_0": value  <=  3;
            "HEIGHT_20_51_1": value  <=  1;
            "HEIGHT_20_52_0": value  <=  4;
            "HEIGHT_20_52_1": value  <=  2;
            "HEIGHT_20_52_2": value  <=  2;
            "HEIGHT_20_53_0": value  <=  7;
            "HEIGHT_20_53_1": value  <=  7;
            "HEIGHT_20_54_0": value  <=  5;
            "HEIGHT_20_54_1": value  <=  5;
            "HEIGHT_20_55_0": value  <=  6;
            "HEIGHT_20_55_1": value  <=  3;
            "HEIGHT_20_55_2": value  <=  3;
            "HEIGHT_20_56_0": value  <=  6;
            "HEIGHT_20_56_1": value  <=  6;
            "HEIGHT_20_57_0": value  <=  2;
            "HEIGHT_20_57_1": value  <=  1;
            "HEIGHT_20_58_0": value  <=  3;
            "HEIGHT_20_58_1": value  <=  3;
            "HEIGHT_20_59_0": value  <=  4;
            "HEIGHT_20_59_1": value  <=  2;
            "HEIGHT_20_60_0": value  <=  1;
            "HEIGHT_20_60_1": value  <=  1;
            "HEIGHT_20_61_0": value  <=  3;
            "HEIGHT_20_61_1": value  <=  1;
            "HEIGHT_20_62_0": value  <=  10;
            "HEIGHT_20_62_1": value  <=  10;
            "HEIGHT_20_63_0": value  <=  6;
            "HEIGHT_20_63_1": value  <=  2;
            "HEIGHT_20_64_0": value  <=  1;
            "HEIGHT_20_64_1": value  <=  1;
            "HEIGHT_20_65_0": value  <=  2;
            "HEIGHT_20_65_1": value  <=  1;
            "HEIGHT_20_66_0": value  <=  2;
            "HEIGHT_20_66_1": value  <=  1;
            "HEIGHT_20_67_0": value  <=  2;
            "HEIGHT_20_67_1": value  <=  1;
            "HEIGHT_20_67_2": value  <=  1;
            "HEIGHT_20_68_0": value  <=  2;
            "HEIGHT_20_68_1": value  <=  1;
            "HEIGHT_20_68_2": value  <=  1;
            "HEIGHT_20_69_0": value  <=  14;
            "HEIGHT_20_69_1": value  <=  14;
            "HEIGHT_20_70_0": value  <=  14;
            "HEIGHT_20_70_1": value  <=  14;
            "HEIGHT_20_71_0": value  <=  14;
            "HEIGHT_20_71_1": value  <=  14;
            "HEIGHT_20_72_0": value  <=  3;
            "HEIGHT_20_72_1": value  <=  1;
            "HEIGHT_20_73_0": value  <=  3;
            "HEIGHT_20_73_1": value  <=  1;
            "HEIGHT_20_74_0": value  <=  16;
            "HEIGHT_20_74_1": value  <=  16;
            "HEIGHT_20_75_0": value  <=  10;
            "HEIGHT_20_75_1": value  <=  5;
            "HEIGHT_20_76_0": value  <=  3;
            "HEIGHT_20_76_1": value  <=  1;
            "HEIGHT_20_77_0": value  <=  12;
            "HEIGHT_20_77_1": value  <=  6;
            "HEIGHT_20_77_2": value  <=  6;
            "HEIGHT_20_78_0": value  <=  2;
            "HEIGHT_20_78_1": value  <=  1;
            "HEIGHT_20_79_0": value  <=  6;
            "HEIGHT_20_79_1": value  <=  3;
            "HEIGHT_20_80_0": value  <=  3;
            "HEIGHT_20_80_1": value  <=  1;
            "HEIGHT_20_81_0": value  <=  6;
            "HEIGHT_20_81_1": value  <=  2;
            "HEIGHT_20_82_0": value  <=  2;
            "HEIGHT_20_82_1": value  <=  1;
            "HEIGHT_20_82_2": value  <=  1;
            "HEIGHT_20_83_0": value  <=  6;
            "HEIGHT_20_83_1": value  <=  2;
            "HEIGHT_20_84_0": value  <=  6;
            "HEIGHT_20_84_1": value  <=  2;
            "HEIGHT_20_85_0": value  <=  6;
            "HEIGHT_20_85_1": value  <=  6;
            "HEIGHT_20_86_0": value  <=  10;
            "HEIGHT_20_86_1": value  <=  5;
            "HEIGHT_20_87_0": value  <=  6;
            "HEIGHT_20_87_1": value  <=  6;
            "HEIGHT_20_88_0": value  <=  3;
            "HEIGHT_20_88_1": value  <=  1;
            "HEIGHT_20_89_0": value  <=  2;
            "HEIGHT_20_89_1": value  <=  1;
            "HEIGHT_20_90_0": value  <=  4;
            "HEIGHT_20_90_1": value  <=  2;
            "HEIGHT_20_90_2": value  <=  2;
            "HEIGHT_20_91_0": value  <=  6;
            "HEIGHT_20_91_1": value  <=  3;
            "HEIGHT_20_91_2": value  <=  3;
            "HEIGHT_20_92_0": value  <=  3;
            "HEIGHT_20_92_1": value  <=  1;
            "HEIGHT_20_93_0": value  <=  3;
            "HEIGHT_20_93_1": value  <=  1;
            "HEIGHT_20_94_0": value  <=  3;
            "HEIGHT_20_94_1": value  <=  1;
            "HEIGHT_20_95_0": value  <=  3;
            "HEIGHT_20_95_1": value  <=  1;
            "HEIGHT_20_96_0": value  <=  4;
            "HEIGHT_20_96_1": value  <=  2;
            "HEIGHT_20_97_0": value  <=  9;
            "HEIGHT_20_97_1": value  <=  3;
            "HEIGHT_20_98_0": value  <=  9;
            "HEIGHT_20_98_1": value  <=  3;
            "HEIGHT_20_99_0": value  <=  1;
            "HEIGHT_20_99_1": value  <=  1;
            "HEIGHT_20_100_0": value  <=  17;
            "HEIGHT_20_100_1": value  <=  17;
            "HEIGHT_20_101_0": value  <=  3;
            "HEIGHT_20_101_1": value  <=  3;
            "HEIGHT_20_102_0": value  <=  4;
            "HEIGHT_20_102_1": value  <=  4;
            "HEIGHT_20_103_0": value  <=  2;
            "HEIGHT_20_103_1": value  <=  1;
            "HEIGHT_20_103_2": value  <=  1;
            "HEIGHT_20_104_0": value  <=  6;
            "HEIGHT_20_104_1": value  <=  2;
            "HEIGHT_20_105_0": value  <=  2;
            "HEIGHT_20_105_1": value  <=  1;
            "HEIGHT_20_106_0": value  <=  14;
            "HEIGHT_20_106_1": value  <=  14;
            "HEIGHT_20_107_0": value  <=  3;
            "HEIGHT_20_107_1": value  <=  1;
            "HEIGHT_20_108_0": value  <=  2;
            "HEIGHT_20_108_1": value  <=  1;
            "HEIGHT_20_109_0": value  <=  8;
            "HEIGHT_20_109_1": value  <=  4;
            "HEIGHT_20_109_2": value  <=  4;
            "HEIGHT_20_110_0": value  <=  3;
            "HEIGHT_20_110_1": value  <=  1;
            "HEIGHT_20_111_0": value  <=  8;
            "HEIGHT_20_111_1": value  <=  4;
            "HEIGHT_20_111_2": value  <=  4;
            "HEIGHT_20_112_0": value  <=  12;
            "HEIGHT_20_112_1": value  <=  6;
            "HEIGHT_20_112_2": value  <=  6;
            "HEIGHT_20_113_0": value  <=  9;
            "HEIGHT_20_113_1": value  <=  3;
            "HEIGHT_20_114_0": value  <=  2;
            "HEIGHT_20_114_1": value  <=  1;
            "HEIGHT_20_115_0": value  <=  6;
            "HEIGHT_20_115_1": value  <=  3;
            "HEIGHT_20_115_2": value  <=  3;
            "HEIGHT_20_116_0": value  <=  2;
            "HEIGHT_20_116_1": value  <=  1;
            "HEIGHT_20_116_2": value  <=  1;
            "HEIGHT_20_117_0": value  <=  6;
            "HEIGHT_20_117_1": value  <=  3;
            "HEIGHT_20_117_2": value  <=  3;
            "HEIGHT_20_118_0": value  <=  2;
            "HEIGHT_20_118_1": value  <=  2;
            "HEIGHT_20_119_0": value  <=  13;
            "HEIGHT_20_119_1": value  <=  13;
            "HEIGHT_20_120_0": value  <=  5;
            "HEIGHT_20_120_1": value  <=  5;
            "HEIGHT_20_121_0": value  <=  10;
            "HEIGHT_20_121_1": value  <=  10;
            "HEIGHT_20_122_0": value  <=  1;
            "HEIGHT_20_122_1": value  <=  1;
            "HEIGHT_20_123_0": value  <=  7;
            "HEIGHT_20_123_1": value  <=  7;
            "HEIGHT_20_124_0": value  <=  7;
            "HEIGHT_20_124_1": value  <=  7;
            "HEIGHT_20_125_0": value  <=  5;
            "HEIGHT_20_125_1": value  <=  5;
            "HEIGHT_20_126_0": value  <=  3;
            "HEIGHT_20_126_1": value  <=  3;
            "HEIGHT_20_127_0": value  <=  6;
            "HEIGHT_20_127_1": value  <=  3;
            "HEIGHT_20_127_2": value  <=  3;
            "HEIGHT_20_128_0": value  <=  4;
            "HEIGHT_20_128_1": value  <=  2;
            "HEIGHT_20_128_2": value  <=  2;
            "HEIGHT_20_129_0": value  <=  2;
            "HEIGHT_20_129_1": value  <=  1;
            "HEIGHT_20_129_2": value  <=  1;
            "HEIGHT_20_130_0": value  <=  12;
            "HEIGHT_20_130_1": value  <=  6;
            "HEIGHT_20_130_2": value  <=  6;
            "HEIGHT_20_131_0": value  <=  3;
            "HEIGHT_20_131_1": value  <=  1;
            "HEIGHT_20_132_0": value  <=  3;
            "HEIGHT_20_132_1": value  <=  1;
            "HEIGHT_20_133_0": value  <=  2;
            "HEIGHT_20_133_1": value  <=  2;
            "HEIGHT_20_134_0": value  <=  2;
            "HEIGHT_20_134_1": value  <=  1;
            "HEIGHT_20_134_2": value  <=  1;
            "HEIGHT_20_135_0": value  <=  3;
            "HEIGHT_20_135_1": value  <=  1;
            "HEIGHT_20_136_0": value  <=  4;
            "HEIGHT_20_136_1": value  <=  2;
            "HEIGHT_20_136_2": value  <=  2;
            "HEIGHT_20_137_0": value  <=  6;
            "HEIGHT_20_137_1": value  <=  3;
            "HEIGHT_20_138_0": value  <=  2;
            "HEIGHT_20_138_1": value  <=  1;
            "HEIGHT_20_139_0": value  <=  6;
            "HEIGHT_20_139_1": value  <=  3;
            "HEIGHT_20_139_2": value  <=  3;
            "HEIGHT_20_140_0": value  <=  4;
            "HEIGHT_20_140_1": value  <=  4;
            "HEIGHT_20_141_0": value  <=  6;
            "HEIGHT_20_141_1": value  <=  3;
            "HEIGHT_20_141_2": value  <=  3;
            "HEIGHT_20_142_0": value  <=  6;
            "HEIGHT_20_142_1": value  <=  2;
            "HEIGHT_20_143_0": value  <=  20;
            "HEIGHT_20_143_1": value  <=  10;
            "HEIGHT_20_144_0": value  <=  6;
            "HEIGHT_20_144_1": value  <=  3;
            "HEIGHT_20_144_2": value  <=  3;
            "HEIGHT_20_145_0": value  <=  6;
            "HEIGHT_20_145_1": value  <=  3;
            "HEIGHT_20_145_2": value  <=  3;
            "HEIGHT_20_146_0": value  <=  1;
            "HEIGHT_20_146_1": value  <=  1;
            "HEIGHT_20_147_0": value  <=  2;
            "HEIGHT_20_147_1": value  <=  2;
            "HEIGHT_20_148_0": value  <=  2;
            "HEIGHT_20_148_1": value  <=  2;
            "HEIGHT_20_149_0": value  <=  6;
            "HEIGHT_20_149_1": value  <=  3;
            "HEIGHT_20_149_2": value  <=  3;
            "HEIGHT_20_150_0": value  <=  6;
            "HEIGHT_20_150_1": value  <=  3;
            "HEIGHT_20_150_2": value  <=  3;
            "HEIGHT_20_151_0": value  <=  6;
            "HEIGHT_20_151_1": value  <=  3;
            "HEIGHT_20_151_2": value  <=  3;
            "HEIGHT_20_152_0": value  <=  6;
            "HEIGHT_20_152_1": value  <=  3;
            "HEIGHT_20_152_2": value  <=  3;
            "HEIGHT_20_153_0": value  <=  12;
            "HEIGHT_20_153_1": value  <=  4;
            "HEIGHT_20_154_0": value  <=  2;
            "HEIGHT_20_154_1": value  <=  2;
            "HEIGHT_20_155_0": value  <=  13;
            "HEIGHT_20_155_1": value  <=  13;
            "HEIGHT_20_156_0": value  <=  13;
            "HEIGHT_20_156_1": value  <=  13;
            "HEIGHT_20_157_0": value  <=  3;
            "HEIGHT_20_157_1": value  <=  1;
            "HEIGHT_20_158_0": value  <=  2;
            "HEIGHT_20_158_1": value  <=  2;
            "HEIGHT_20_159_0": value  <=  8;
            "HEIGHT_20_159_1": value  <=  4;
            "HEIGHT_20_159_2": value  <=  4;
            "HEIGHT_20_160_0": value  <=  5;
            "HEIGHT_20_160_1": value  <=  5;
            "HEIGHT_20_161_0": value  <=  7;
            "HEIGHT_20_161_1": value  <=  7;
            "HEIGHT_20_162_0": value  <=  2;
            "HEIGHT_20_162_1": value  <=  2;
            "HEIGHT_20_163_0": value  <=  3;
            "HEIGHT_20_163_1": value  <=  1;
            "HEIGHT_20_164_0": value  <=  3;
            "HEIGHT_20_164_1": value  <=  1;
            "HEIGHT_20_165_0": value  <=  3;
            "HEIGHT_20_165_1": value  <=  1;
            "HEIGHT_20_166_0": value  <=  12;
            "HEIGHT_20_166_1": value  <=  4;
            "HEIGHT_20_167_0": value  <=  3;
            "HEIGHT_20_167_1": value  <=  1;
            "HEIGHT_20_168_0": value  <=  3;
            "HEIGHT_20_168_1": value  <=  1;
            "HEIGHT_20_169_0": value  <=  3;
            "HEIGHT_20_169_1": value  <=  1;
            "HEIGHT_20_170_0": value  <=  7;
            "HEIGHT_20_170_1": value  <=  7;
            "HEIGHT_20_171_0": value  <=  8;
            "HEIGHT_20_171_1": value  <=  4;
            "HEIGHT_20_171_2": value  <=  4;
            "HEIGHT_20_172_0": value  <=  3;
            "HEIGHT_20_172_1": value  <=  1;
            "HEIGHT_20_173_0": value  <=  2;
            "HEIGHT_20_173_1": value  <=  1;
            "HEIGHT_20_173_2": value  <=  1;
            "HEIGHT_20_174_0": value  <=  3;
            "HEIGHT_20_174_1": value  <=  1;
            "HEIGHT_20_175_0": value  <=  3;
            "HEIGHT_20_175_1": value  <=  3;
            "HEIGHT_20_176_0": value  <=  3;
            "HEIGHT_20_176_1": value  <=  1;
            "HEIGHT_20_177_0": value  <=  3;
            "HEIGHT_20_177_1": value  <=  1;
            "HEIGHT_20_178_0": value  <=  3;
            "HEIGHT_20_178_1": value  <=  1;
            "HEIGHT_20_179_0": value  <=  8;
            "HEIGHT_20_179_1": value  <=  4;
            "HEIGHT_20_179_2": value  <=  4;
            "HEIGHT_20_180_0": value  <=  8;
            "HEIGHT_20_180_1": value  <=  4;
            "HEIGHT_20_180_2": value  <=  4;
            "HEIGHT_20_181_0": value  <=  6;
            "HEIGHT_20_181_1": value  <=  2;
            "HEIGHT_20_182_0": value  <=  6;
            "HEIGHT_20_182_1": value  <=  2;
            "HEIGHT_20_183_0": value  <=  2;
            "HEIGHT_20_183_1": value  <=  1;
            "HEIGHT_20_183_2": value  <=  1;
            "HEIGHT_20_184_0": value  <=  6;
            "HEIGHT_20_184_1": value  <=  3;
            "HEIGHT_20_185_0": value  <=  3;
            "HEIGHT_20_185_1": value  <=  1;
            "HEIGHT_20_186_0": value  <=  2;
            "HEIGHT_20_186_1": value  <=  1;
            "HEIGHT_20_186_2": value  <=  1;
            "HEIGHT_20_187_0": value  <=  3;
            "HEIGHT_20_187_1": value  <=  1;
            "HEIGHT_20_188_0": value  <=  2;
            "HEIGHT_20_188_1": value  <=  1;
            "HEIGHT_20_188_2": value  <=  1;
            "HEIGHT_20_189_0": value  <=  3;
            "HEIGHT_20_189_1": value  <=  1;
            "HEIGHT_20_190_0": value  <=  2;
            "HEIGHT_20_190_1": value  <=  2;
            "HEIGHT_20_191_0": value  <=  3;
            "HEIGHT_20_191_1": value  <=  3;
            "HEIGHT_20_192_0": value  <=  2;
            "HEIGHT_20_192_1": value  <=  1;
            "HEIGHT_20_192_2": value  <=  1;
            "HEIGHT_20_193_0": value  <=  4;
            "HEIGHT_20_193_1": value  <=  4;
            "HEIGHT_20_194_0": value  <=  3;
            "HEIGHT_20_194_1": value  <=  1;
            "HEIGHT_20_195_0": value  <=  2;
            "HEIGHT_20_195_1": value  <=  1;
            "HEIGHT_20_196_0": value  <=  2;
            "HEIGHT_20_196_1": value  <=  1;
            "HEIGHT_20_196_2": value  <=  1;
            "HEIGHT_20_197_0": value  <=  4;
            "HEIGHT_20_197_1": value  <=  4;
            "HEIGHT_20_198_0": value  <=  6;
            "HEIGHT_20_198_1": value  <=  6;
            "HEIGHT_20_199_0": value  <=  2;
            "HEIGHT_20_199_1": value  <=  1;
            "HEIGHT_20_200_0": value  <=  4;
            "HEIGHT_20_200_1": value  <=  2;
            "HEIGHT_20_200_2": value  <=  2;
            "HEIGHT_20_201_0": value  <=  2;
            "HEIGHT_20_201_1": value  <=  1;
            "HEIGHT_20_201_2": value  <=  1;
            "HEIGHT_20_202_0": value  <=  2;
            "HEIGHT_20_202_1": value  <=  1;
            "HEIGHT_20_203_0": value  <=  14;
            "HEIGHT_20_203_1": value  <=  14;
            "HEIGHT_20_204_0": value  <=  3;
            "HEIGHT_20_204_1": value  <=  1;
            "HEIGHT_20_205_0": value  <=  14;
            "HEIGHT_20_205_1": value  <=  14;
            "HEIGHT_20_206_0": value  <=  7;
            "HEIGHT_20_206_1": value  <=  7;
            "HEIGHT_20_207_0": value  <=  2;
            "HEIGHT_20_207_1": value  <=  1;
            "HEIGHT_20_208_0": value  <=  1;
            "HEIGHT_20_208_1": value  <=  1;
            "HEIGHT_20_209_0": value  <=  4;
            "HEIGHT_20_209_1": value  <=  4;
            "HEIGHT_20_210_0": value  <=  2;
            "HEIGHT_20_210_1": value  <=  1;
            "HEIGHT_21_0_0": value  <=  9;
            "HEIGHT_21_0_1": value  <=  3;
            "HEIGHT_21_1_0": value  <=  10;
            "HEIGHT_21_1_1": value  <=  10;
            "HEIGHT_21_2_0": value  <=  7;
            "HEIGHT_21_2_1": value  <=  7;
            "HEIGHT_21_3_0": value  <=  1;
            "HEIGHT_21_3_1": value  <=  1;
            "HEIGHT_21_4_0": value  <=  1;
            "HEIGHT_21_4_1": value  <=  1;
            "HEIGHT_21_5_0": value  <=  4;
            "HEIGHT_21_5_1": value  <=  2;
            "HEIGHT_21_6_0": value  <=  4;
            "HEIGHT_21_6_1": value  <=  4;
            "HEIGHT_21_7_0": value  <=  6;
            "HEIGHT_21_7_1": value  <=  3;
            "HEIGHT_21_8_0": value  <=  3;
            "HEIGHT_21_8_1": value  <=  1;
            "HEIGHT_21_9_0": value  <=  16;
            "HEIGHT_21_9_1": value  <=  8;
            "HEIGHT_21_9_2": value  <=  8;
            "HEIGHT_21_10_0": value  <=  6;
            "HEIGHT_21_10_1": value  <=  3;
            "HEIGHT_21_11_0": value  <=  2;
            "HEIGHT_21_11_1": value  <=  1;
            "HEIGHT_21_12_0": value  <=  2;
            "HEIGHT_21_12_1": value  <=  1;
            "HEIGHT_21_12_2": value  <=  1;
            "HEIGHT_21_13_0": value  <=  10;
            "HEIGHT_21_13_1": value  <=  5;
            "HEIGHT_21_13_2": value  <=  5;
            "HEIGHT_21_14_0": value  <=  10;
            "HEIGHT_21_14_1": value  <=  5;
            "HEIGHT_21_15_0": value  <=  2;
            "HEIGHT_21_15_1": value  <=  2;
            "HEIGHT_21_16_0": value  <=  2;
            "HEIGHT_21_16_1": value  <=  2;
            "HEIGHT_21_17_0": value  <=  6;
            "HEIGHT_21_17_1": value  <=  2;
            "HEIGHT_21_18_0": value  <=  2;
            "HEIGHT_21_18_1": value  <=  2;
            "HEIGHT_21_19_0": value  <=  3;
            "HEIGHT_21_19_1": value  <=  1;
            "HEIGHT_21_20_0": value  <=  3;
            "HEIGHT_21_20_1": value  <=  1;
            "HEIGHT_21_21_0": value  <=  2;
            "HEIGHT_21_21_1": value  <=  1;
            "HEIGHT_21_22_0": value  <=  18;
            "HEIGHT_21_22_1": value  <=  6;
            "HEIGHT_21_23_0": value  <=  2;
            "HEIGHT_21_23_1": value  <=  2;
            "HEIGHT_21_24_0": value  <=  3;
            "HEIGHT_21_24_1": value  <=  1;
            "HEIGHT_21_25_0": value  <=  6;
            "HEIGHT_21_25_1": value  <=  2;
            "HEIGHT_21_26_0": value  <=  4;
            "HEIGHT_21_26_1": value  <=  4;
            "HEIGHT_21_27_0": value  <=  2;
            "HEIGHT_21_27_1": value  <=  1;
            "HEIGHT_21_28_0": value  <=  2;
            "HEIGHT_21_28_1": value  <=  1;
            "HEIGHT_21_29_0": value  <=  3;
            "HEIGHT_21_29_1": value  <=  1;
            "HEIGHT_21_30_0": value  <=  3;
            "HEIGHT_21_30_1": value  <=  1;
            "HEIGHT_21_31_0": value  <=  3;
            "HEIGHT_21_31_1": value  <=  1;
            "HEIGHT_21_32_0": value  <=  3;
            "HEIGHT_21_32_1": value  <=  1;
            "HEIGHT_21_33_0": value  <=  4;
            "HEIGHT_21_33_1": value  <=  2;
            "HEIGHT_21_33_2": value  <=  2;
            "HEIGHT_21_34_0": value  <=  6;
            "HEIGHT_21_34_1": value  <=  3;
            "HEIGHT_21_35_0": value  <=  2;
            "HEIGHT_21_35_1": value  <=  1;
            "HEIGHT_21_35_2": value  <=  1;
            "HEIGHT_21_36_0": value  <=  3;
            "HEIGHT_21_36_1": value  <=  1;
            "HEIGHT_21_37_0": value  <=  6;
            "HEIGHT_21_37_1": value  <=  2;
            "HEIGHT_21_38_0": value  <=  3;
            "HEIGHT_21_38_1": value  <=  1;
            "HEIGHT_21_39_0": value  <=  6;
            "HEIGHT_21_39_1": value  <=  2;
            "HEIGHT_21_40_0": value  <=  6;
            "HEIGHT_21_40_1": value  <=  2;
            "HEIGHT_21_41_0": value  <=  3;
            "HEIGHT_21_41_1": value  <=  3;
            "HEIGHT_21_42_0": value  <=  1;
            "HEIGHT_21_42_1": value  <=  1;
            "HEIGHT_21_43_0": value  <=  3;
            "HEIGHT_21_43_1": value  <=  1;
            "HEIGHT_21_44_0": value  <=  6;
            "HEIGHT_21_44_1": value  <=  2;
            "HEIGHT_21_45_0": value  <=  2;
            "HEIGHT_21_45_1": value  <=  1;
            "HEIGHT_21_46_0": value  <=  2;
            "HEIGHT_21_46_1": value  <=  1;
            "HEIGHT_21_47_0": value  <=  8;
            "HEIGHT_21_47_1": value  <=  4;
            "HEIGHT_21_47_2": value  <=  4;
            "HEIGHT_21_48_0": value  <=  6;
            "HEIGHT_21_48_1": value  <=  3;
            "HEIGHT_21_48_2": value  <=  3;
            "HEIGHT_21_49_0": value  <=  1;
            "HEIGHT_21_49_1": value  <=  1;
            "HEIGHT_21_50_0": value  <=  10;
            "HEIGHT_21_50_1": value  <=  5;
            "HEIGHT_21_50_2": value  <=  5;
            "HEIGHT_21_51_0": value  <=  6;
            "HEIGHT_21_51_1": value  <=  6;
            "HEIGHT_21_52_0": value  <=  6;
            "HEIGHT_21_52_1": value  <=  2;
            "HEIGHT_21_53_0": value  <=  2;
            "HEIGHT_21_53_1": value  <=  1;
            "HEIGHT_21_54_0": value  <=  6;
            "HEIGHT_21_54_1": value  <=  3;
            "HEIGHT_21_54_2": value  <=  3;
            "HEIGHT_21_55_0": value  <=  6;
            "HEIGHT_21_55_1": value  <=  6;
            "HEIGHT_21_56_0": value  <=  2;
            "HEIGHT_21_56_1": value  <=  1;
            "HEIGHT_21_57_0": value  <=  3;
            "HEIGHT_21_57_1": value  <=  3;
            "HEIGHT_21_58_0": value  <=  3;
            "HEIGHT_21_58_1": value  <=  1;
            "HEIGHT_21_59_0": value  <=  3;
            "HEIGHT_21_59_1": value  <=  3;
            "HEIGHT_21_60_0": value  <=  9;
            "HEIGHT_21_60_1": value  <=  9;
            "HEIGHT_21_61_0": value  <=  15;
            "HEIGHT_21_61_1": value  <=  15;
            "HEIGHT_21_62_0": value  <=  15;
            "HEIGHT_21_62_1": value  <=  15;
            "HEIGHT_21_63_0": value  <=  3;
            "HEIGHT_21_63_1": value  <=  3;
            "HEIGHT_21_64_0": value  <=  3;
            "HEIGHT_21_64_1": value  <=  3;
            "HEIGHT_21_65_0": value  <=  2;
            "HEIGHT_21_65_1": value  <=  1;
            "HEIGHT_21_65_2": value  <=  1;
            "HEIGHT_21_66_0": value  <=  2;
            "HEIGHT_21_66_1": value  <=  1;
            "HEIGHT_21_66_2": value  <=  1;
            "HEIGHT_21_67_0": value  <=  4;
            "HEIGHT_21_67_1": value  <=  4;
            "HEIGHT_21_68_0": value  <=  3;
            "HEIGHT_21_68_1": value  <=  1;
            "HEIGHT_21_69_0": value  <=  2;
            "HEIGHT_21_69_1": value  <=  1;
            "HEIGHT_21_70_0": value  <=  2;
            "HEIGHT_21_70_1": value  <=  2;
            "HEIGHT_21_71_0": value  <=  2;
            "HEIGHT_21_71_1": value  <=  2;
            "HEIGHT_21_72_0": value  <=  2;
            "HEIGHT_21_72_1": value  <=  2;
            "HEIGHT_21_73_0": value  <=  4;
            "HEIGHT_21_73_1": value  <=  4;
            "HEIGHT_21_74_0": value  <=  4;
            "HEIGHT_21_74_1": value  <=  4;
            "HEIGHT_21_75_0": value  <=  4;
            "HEIGHT_21_75_1": value  <=  2;
            "HEIGHT_21_75_2": value  <=  2;
            "HEIGHT_21_76_0": value  <=  3;
            "HEIGHT_21_76_1": value  <=  1;
            "HEIGHT_21_77_0": value  <=  8;
            "HEIGHT_21_77_1": value  <=  4;
            "HEIGHT_21_78_0": value  <=  8;
            "HEIGHT_21_78_1": value  <=  4;
            "HEIGHT_21_78_2": value  <=  4;
            "HEIGHT_21_79_0": value  <=  1;
            "HEIGHT_21_79_1": value  <=  1;
            "HEIGHT_21_80_0": value  <=  6;
            "HEIGHT_21_80_1": value  <=  3;
            "HEIGHT_21_81_0": value  <=  1;
            "HEIGHT_21_81_1": value  <=  1;
            "HEIGHT_21_82_0": value  <=  1;
            "HEIGHT_21_82_1": value  <=  1;
            "HEIGHT_21_83_0": value  <=  14;
            "HEIGHT_21_83_1": value  <=  7;
            "HEIGHT_21_84_0": value  <=  10;
            "HEIGHT_21_84_1": value  <=  5;
            "HEIGHT_21_84_2": value  <=  5;
            "HEIGHT_21_85_0": value  <=  3;
            "HEIGHT_21_85_1": value  <=  1;
            "HEIGHT_21_86_0": value  <=  3;
            "HEIGHT_21_86_1": value  <=  3;
            "HEIGHT_21_87_0": value  <=  3;
            "HEIGHT_21_87_1": value  <=  1;
            "HEIGHT_21_88_0": value  <=  3;
            "HEIGHT_21_88_1": value  <=  1;
            "HEIGHT_21_89_0": value  <=  2;
            "HEIGHT_21_89_1": value  <=  1;
            "HEIGHT_21_89_2": value  <=  1;
            "HEIGHT_21_90_0": value  <=  1;
            "HEIGHT_21_90_1": value  <=  1;
            "HEIGHT_21_91_0": value  <=  4;
            "HEIGHT_21_91_1": value  <=  2;
            "HEIGHT_21_92_0": value  <=  3;
            "HEIGHT_21_92_1": value  <=  1;
            "HEIGHT_21_93_0": value  <=  4;
            "HEIGHT_21_93_1": value  <=  4;
            "HEIGHT_21_94_0": value  <=  10;
            "HEIGHT_21_94_1": value  <=  10;
            "HEIGHT_21_95_0": value  <=  4;
            "HEIGHT_21_95_1": value  <=  4;
            "HEIGHT_21_96_0": value  <=  4;
            "HEIGHT_21_96_1": value  <=  4;
            "HEIGHT_21_97_0": value  <=  3;
            "HEIGHT_21_97_1": value  <=  3;
            "HEIGHT_21_98_0": value  <=  3;
            "HEIGHT_21_98_1": value  <=  3;
            "HEIGHT_21_99_0": value  <=  2;
            "HEIGHT_21_99_1": value  <=  2;
            "HEIGHT_21_100_0": value  <=  2;
            "HEIGHT_21_100_1": value  <=  2;
            "HEIGHT_21_101_0": value  <=  2;
            "HEIGHT_21_101_1": value  <=  1;
            "HEIGHT_21_102_0": value  <=  6;
            "HEIGHT_21_102_1": value  <=  3;
            "HEIGHT_21_102_2": value  <=  3;
            "HEIGHT_21_103_0": value  <=  2;
            "HEIGHT_21_103_1": value  <=  1;
            "HEIGHT_21_103_2": value  <=  1;
            "HEIGHT_21_104_0": value  <=  3;
            "HEIGHT_21_104_1": value  <=  1;
            "HEIGHT_21_105_0": value  <=  2;
            "HEIGHT_21_105_1": value  <=  2;
            "HEIGHT_21_106_0": value  <=  12;
            "HEIGHT_21_106_1": value  <=  6;
            "HEIGHT_21_107_0": value  <=  2;
            "HEIGHT_21_107_1": value  <=  1;
            "HEIGHT_21_108_0": value  <=  2;
            "HEIGHT_21_108_1": value  <=  1;
            "HEIGHT_21_109_0": value  <=  3;
            "HEIGHT_21_109_1": value  <=  1;
            "HEIGHT_21_110_0": value  <=  3;
            "HEIGHT_21_110_1": value  <=  1;
            "HEIGHT_21_111_0": value  <=  3;
            "HEIGHT_21_111_1": value  <=  1;
            "HEIGHT_21_112_0": value  <=  3;
            "HEIGHT_21_112_1": value  <=  1;
            "HEIGHT_21_113_0": value  <=  6;
            "HEIGHT_21_113_1": value  <=  3;
            "HEIGHT_21_113_2": value  <=  3;
            "HEIGHT_21_114_0": value  <=  2;
            "HEIGHT_21_114_1": value  <=  2;
            "HEIGHT_21_115_0": value  <=  6;
            "HEIGHT_21_115_1": value  <=  6;
            "HEIGHT_21_116_0": value  <=  6;
            "HEIGHT_21_116_1": value  <=  6;
            "HEIGHT_21_117_0": value  <=  2;
            "HEIGHT_21_117_1": value  <=  1;
            "HEIGHT_21_118_0": value  <=  2;
            "HEIGHT_21_118_1": value  <=  1;
            "HEIGHT_21_119_0": value  <=  2;
            "HEIGHT_21_119_1": value  <=  1;
            "HEIGHT_21_120_0": value  <=  2;
            "HEIGHT_21_120_1": value  <=  1;
            "HEIGHT_21_120_2": value  <=  1;
            "HEIGHT_21_121_0": value  <=  7;
            "HEIGHT_21_121_1": value  <=  7;
            "HEIGHT_21_122_0": value  <=  2;
            "HEIGHT_21_122_1": value  <=  1;
            "HEIGHT_21_123_0": value  <=  7;
            "HEIGHT_21_123_1": value  <=  7;
            "HEIGHT_21_124_0": value  <=  16;
            "HEIGHT_21_124_1": value  <=  8;
            "HEIGHT_21_124_2": value  <=  8;
            "HEIGHT_21_125_0": value  <=  7;
            "HEIGHT_21_125_1": value  <=  7;
            "HEIGHT_21_126_0": value  <=  7;
            "HEIGHT_21_126_1": value  <=  7;
            "HEIGHT_21_127_0": value  <=  4;
            "HEIGHT_21_127_1": value  <=  4;
            "HEIGHT_21_128_0": value  <=  4;
            "HEIGHT_21_128_1": value  <=  4;
            "HEIGHT_21_129_0": value  <=  7;
            "HEIGHT_21_129_1": value  <=  7;
            "HEIGHT_21_130_0": value  <=  7;
            "HEIGHT_21_130_1": value  <=  7;
            "HEIGHT_21_131_0": value  <=  14;
            "HEIGHT_21_131_1": value  <=  7;
            "HEIGHT_21_132_0": value  <=  4;
            "HEIGHT_21_132_1": value  <=  2;
            "HEIGHT_21_133_0": value  <=  2;
            "HEIGHT_21_133_1": value  <=  1;
            "HEIGHT_21_134_0": value  <=  6;
            "HEIGHT_21_134_1": value  <=  3;
            "HEIGHT_21_134_2": value  <=  3;
            "HEIGHT_21_135_0": value  <=  2;
            "HEIGHT_21_135_1": value  <=  1;
            "HEIGHT_21_136_0": value  <=  14;
            "HEIGHT_21_136_1": value  <=  7;
            "HEIGHT_21_137_0": value  <=  12;
            "HEIGHT_21_137_1": value  <=  12;
            "HEIGHT_21_138_0": value  <=  3;
            "HEIGHT_21_138_1": value  <=  1;
            "HEIGHT_21_139_0": value  <=  16;
            "HEIGHT_21_139_1": value  <=  8;
            "HEIGHT_21_140_0": value  <=  12;
            "HEIGHT_21_140_1": value  <=  12;
            "HEIGHT_21_141_0": value  <=  7;
            "HEIGHT_21_141_1": value  <=  7;
            "HEIGHT_21_142_0": value  <=  2;
            "HEIGHT_21_142_1": value  <=  1;
            "HEIGHT_21_143_0": value  <=  6;
            "HEIGHT_21_143_1": value  <=  2;
            "HEIGHT_21_144_0": value  <=  2;
            "HEIGHT_21_144_1": value  <=  1;
            "HEIGHT_21_145_0": value  <=  9;
            "HEIGHT_21_145_1": value  <=  3;
            "HEIGHT_21_146_0": value  <=  1;
            "HEIGHT_21_146_1": value  <=  1;
            "HEIGHT_21_147_0": value  <=  4;
            "HEIGHT_21_147_1": value  <=  2;
            "HEIGHT_21_147_2": value  <=  2;
            "HEIGHT_21_148_0": value  <=  12;
            "HEIGHT_21_148_1": value  <=  4;
            "HEIGHT_21_149_0": value  <=  12;
            "HEIGHT_21_149_1": value  <=  4;
            "HEIGHT_21_150_0": value  <=  3;
            "HEIGHT_21_150_1": value  <=  1;
            "HEIGHT_21_151_0": value  <=  3;
            "HEIGHT_21_151_1": value  <=  1;
            "HEIGHT_21_152_0": value  <=  3;
            "HEIGHT_21_152_1": value  <=  1;
            "HEIGHT_21_153_0": value  <=  6;
            "HEIGHT_21_153_1": value  <=  2;
            "HEIGHT_21_154_0": value  <=  6;
            "HEIGHT_21_154_1": value  <=  2;
            "HEIGHT_21_155_0": value  <=  3;
            "HEIGHT_21_155_1": value  <=  1;
            "HEIGHT_21_156_0": value  <=  3;
            "HEIGHT_21_156_1": value  <=  1;
            "HEIGHT_21_157_0": value  <=  6;
            "HEIGHT_21_157_1": value  <=  2;
            "HEIGHT_21_158_0": value  <=  9;
            "HEIGHT_21_158_1": value  <=  9;
            "HEIGHT_21_159_0": value  <=  2;
            "HEIGHT_21_159_1": value  <=  2;
            "HEIGHT_21_160_0": value  <=  2;
            "HEIGHT_21_160_1": value  <=  1;
            "HEIGHT_21_160_2": value  <=  1;
            "HEIGHT_21_161_0": value  <=  3;
            "HEIGHT_21_161_1": value  <=  1;
            "HEIGHT_21_162_0": value  <=  3;
            "HEIGHT_21_162_1": value  <=  1;
            "HEIGHT_21_163_0": value  <=  2;
            "HEIGHT_21_163_1": value  <=  1;
            "HEIGHT_21_164_0": value  <=  3;
            "HEIGHT_21_164_1": value  <=  1;
            "HEIGHT_21_165_0": value  <=  6;
            "HEIGHT_21_165_1": value  <=  3;
            "HEIGHT_21_166_0": value  <=  4;
            "HEIGHT_21_166_1": value  <=  2;
            "HEIGHT_21_166_2": value  <=  2;
            "HEIGHT_21_167_0": value  <=  7;
            "HEIGHT_21_167_1": value  <=  7;
            "HEIGHT_21_168_0": value  <=  2;
            "HEIGHT_21_168_1": value  <=  1;
            "HEIGHT_21_169_0": value  <=  10;
            "HEIGHT_21_169_1": value  <=  5;
            "HEIGHT_21_170_0": value  <=  2;
            "HEIGHT_21_170_1": value  <=  1;
            "HEIGHT_21_171_0": value  <=  9;
            "HEIGHT_21_171_1": value  <=  3;
            "HEIGHT_21_172_0": value  <=  7;
            "HEIGHT_21_172_1": value  <=  7;
            "HEIGHT_21_173_0": value  <=  12;
            "HEIGHT_21_173_1": value  <=  6;
            "HEIGHT_21_173_2": value  <=  6;
            "HEIGHT_21_174_0": value  <=  4;
            "HEIGHT_21_174_1": value  <=  2;
            "HEIGHT_21_175_0": value  <=  3;
            "HEIGHT_21_175_1": value  <=  1;
            "HEIGHT_21_176_0": value  <=  7;
            "HEIGHT_21_176_1": value  <=  7;
            "HEIGHT_21_177_0": value  <=  4;
            "HEIGHT_21_177_1": value  <=  4;
            "HEIGHT_21_178_0": value  <=  4;
            "HEIGHT_21_178_1": value  <=  4;
            "HEIGHT_21_179_0": value  <=  1;
            "HEIGHT_21_179_1": value  <=  1;
            "HEIGHT_21_180_0": value  <=  4;
            "HEIGHT_21_180_1": value  <=  2;
            "HEIGHT_21_180_2": value  <=  2;
            "HEIGHT_21_181_0": value  <=  6;
            "HEIGHT_21_181_1": value  <=  3;
            "HEIGHT_21_181_2": value  <=  3;
            "HEIGHT_21_182_0": value  <=  8;
            "HEIGHT_21_182_1": value  <=  4;
            "HEIGHT_21_183_0": value  <=  8;
            "HEIGHT_21_183_1": value  <=  4;
            "HEIGHT_21_183_2": value  <=  4;
            "HEIGHT_21_184_0": value  <=  8;
            "HEIGHT_21_184_1": value  <=  4;
            "HEIGHT_21_184_2": value  <=  4;
            "HEIGHT_21_185_0": value  <=  3;
            "HEIGHT_21_185_1": value  <=  1;
            "HEIGHT_21_186_0": value  <=  10;
            "HEIGHT_21_186_1": value  <=  5;
            "HEIGHT_21_187_0": value  <=  2;
            "HEIGHT_21_187_1": value  <=  1;
            "HEIGHT_21_188_0": value  <=  8;
            "HEIGHT_21_188_1": value  <=  4;
            "HEIGHT_21_189_0": value  <=  6;
            "HEIGHT_21_189_1": value  <=  3;
            "HEIGHT_21_190_0": value  <=  3;
            "HEIGHT_21_190_1": value  <=  1;
            "HEIGHT_21_191_0": value  <=  2;
            "HEIGHT_21_191_1": value  <=  1;
            "HEIGHT_21_192_0": value  <=  2;
            "HEIGHT_21_192_1": value  <=  2;
            "HEIGHT_21_193_0": value  <=  14;
            "HEIGHT_21_193_1": value  <=  7;
            "HEIGHT_21_194_0": value  <=  1;
            "HEIGHT_21_194_1": value  <=  1;
            "HEIGHT_21_195_0": value  <=  2;
            "HEIGHT_21_195_1": value  <=  2;
            "HEIGHT_21_196_0": value  <=  9;
            "HEIGHT_21_196_1": value  <=  9;
            "HEIGHT_21_197_0": value  <=  3;
            "HEIGHT_21_197_1": value  <=  1;
            "HEIGHT_21_198_0": value  <=  1;
            "HEIGHT_21_198_1": value  <=  1;
            "HEIGHT_21_199_0": value  <=  4;
            "HEIGHT_21_199_1": value  <=  4;
            "HEIGHT_21_200_0": value  <=  6;
            "HEIGHT_21_200_1": value  <=  6;
            "HEIGHT_21_201_0": value  <=  4;
            "HEIGHT_21_201_1": value  <=  4;
            "HEIGHT_21_202_0": value  <=  4;
            "HEIGHT_21_202_1": value  <=  4;
            "HEIGHT_21_203_0": value  <=  9;
            "HEIGHT_21_203_1": value  <=  3;
            "HEIGHT_21_204_0": value  <=  3;
            "HEIGHT_21_204_1": value  <=  1;
            "HEIGHT_21_205_0": value  <=  2;
            "HEIGHT_21_205_1": value  <=  1;
            "HEIGHT_21_206_0": value  <=  3;
            "HEIGHT_21_206_1": value  <=  3;
            "HEIGHT_21_207_0": value  <=  6;
            "HEIGHT_21_207_1": value  <=  6;
            "HEIGHT_21_208_0": value  <=  3;
            "HEIGHT_21_208_1": value  <=  1;
            "HEIGHT_21_209_0": value  <=  3;
            "HEIGHT_21_209_1": value  <=  1;
            "HEIGHT_21_210_0": value  <=  4;
            "HEIGHT_21_210_1": value  <=  2;
            "HEIGHT_21_211_0": value  <=  6;
            "HEIGHT_21_211_1": value  <=  3;
            "HEIGHT_21_212_0": value  <=  6;
            "HEIGHT_21_212_1": value  <=  3;
            "HEIGHT_21_212_2": value  <=  3;

            default: value <= -1;

        endcase

    end

endmodule 
