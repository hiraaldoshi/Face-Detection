module Right (

input string name,
output real value

);

always_comb
    begin

        case (name)

            RIGHT_0_0: value  <= 0.83781069517135620117;
            RIGHT_0_1: value  <= 0.74888122081756591797;
            RIGHT_0_2: value  <= 0.63748198747634887695;
            RIGHT_1_0: value  <= 0.71109461784362792969;
            RIGHT_1_1: value  <= 0.66686922311782836914;
            RIGHT_1_2: value  <= 0.65540069341659545898;
            RIGHT_1_3: value  <= 0.09141451865434649382;
            RIGHT_1_4: value  <= 0.60318958759307861328;
            RIGHT_1_5: value  <= 0.79203182458877563477;
            RIGHT_1_6: value  <= 0.20885099470615389738;
            RIGHT_1_7: value  <= 0.63602739572525024414;
            RIGHT_1_8: value  <= 0.58007007837295532227;
            RIGHT_1_9: value  <= 0.57870548963546752930;
            RIGHT_1_10: value  <= 0.13622370362281799316;
            RIGHT_1_11: value  <= 0.47177401185035711118;
            RIGHT_1_12: value  <= 0.28345298767089838199;
            RIGHT_1_13: value  <= 0.70600342750549316406;
            RIGHT_1_14: value  <= 0.60515749454498291016;
            RIGHT_1_15: value  <= 0.56752568483352661133;
            RIGHT_2_0: value  <= 0.14248579740524289217;
            RIGHT_2_1: value  <= 0.12884770333766940031;
            RIGHT_2_2: value  <= 0.61931931972503662109;
            RIGHT_2_3: value  <= 0.56700158119201660156;
            RIGHT_2_4: value  <= 0.59052079916000366211;
            RIGHT_2_5: value  <= 0.57388240098953247070;
            RIGHT_2_6: value  <= 0.57827740907669067383;
            RIGHT_2_7: value  <= 0.56954258680343627930;
            RIGHT_2_8: value  <= 0.59566420316696166992;
            RIGHT_2_9: value  <= 0.55220472812652587891;
            RIGHT_2_10: value  <= 0.55590140819549560547;
            RIGHT_2_11: value  <= 0.61888492107391357422;
            RIGHT_2_12: value  <= 0.54759448766708374023;
            RIGHT_2_13: value  <= 0.57113999128341674805;
            RIGHT_2_14: value  <= 0.33180978894233698062;
            RIGHT_2_15: value  <= 0.56028461456298828125;
            RIGHT_2_16: value  <= 0.61317151784896850586;
            RIGHT_2_17: value  <= 0.34595629572868352719;
            RIGHT_2_18: value  <= 0.69908452033996582031;
            RIGHT_2_19: value  <= 0.78014570474624633789;
            RIGHT_2_20: value  <= 0.13198269903659820557;
            RIGHT_3_0: value  <= 0.61998707056045532227;
            RIGHT_3_1: value  <= 0.18849289417266851254;
            RIGHT_3_2: value  <= 0.58579277992248535156;
            RIGHT_3_3: value  <= 0.63592398166656494141;
            RIGHT_3_4: value  <= 0.21756289899349209871;
            RIGHT_3_5: value  <= 0.29795908927917480469;
            RIGHT_3_6: value  <= 0.58766472339630126953;
            RIGHT_3_7: value  <= 0.51942020654678344727;
            RIGHT_3_8: value  <= 0.58174091577529907227;
            RIGHT_3_9: value  <= 0.56985449790954589844;
            RIGHT_3_10: value  <= 0.75593662261962890625;
            RIGHT_3_11: value  <= 0.56134271621704101562;
            RIGHT_3_12: value  <= 0.26427671313285827637;
            RIGHT_3_13: value  <= 0.27517059445381170102;
            RIGHT_3_14: value  <= 0.57525688409805297852;
            RIGHT_3_15: value  <= 0.23348769545555120297;
            RIGHT_3_16: value  <= 0.20631550252437588777;
            RIGHT_3_17: value  <= 0.30688610672950750180;
            RIGHT_3_18: value  <= 0.61128681898117065430;
            RIGHT_3_19: value  <= 0.60252362489700317383;
            RIGHT_3_20: value  <= 0.53628271818161010742;
            RIGHT_3_21: value  <= 0.55293101072311401367;
            RIGHT_3_22: value  <= 0.71018958091735839844;
            RIGHT_3_23: value  <= 0.63919639587402343750;
            RIGHT_3_24: value  <= 0.54337137937545776367;
            RIGHT_3_25: value  <= 0.32391890883445739746;
            RIGHT_3_26: value  <= 0.29118689894676208496;
            RIGHT_3_27: value  <= 0.51966291666030883789;
            RIGHT_3_28: value  <= 0.55335938930511474609;
            RIGHT_3_29: value  <= 0.69753772020339965820;
            RIGHT_3_30: value  <= 0.54979521036148071289;
            RIGHT_3_31: value  <= 0.23855470120906829834;
            RIGHT_3_32: value  <= 0.69836008548736572266;
            RIGHT_3_33: value  <= 0.53909200429916381836;
            RIGHT_3_34: value  <= 0.31203660368919372559;
            RIGHT_3_35: value  <= 0.17706030607223510742;
            RIGHT_3_36: value  <= 0.12110190093517300691;
            RIGHT_3_37: value  <= 0.33112218976020807437;
            RIGHT_3_38: value  <= 0.44519689679145807437;
            RIGHT_4_0: value  <= 0.60767322778701782227;
            RIGHT_4_1: value  <= 0.12553839385509490967;
            RIGHT_4_2: value  <= 0.57289612293243408203;
            RIGHT_4_3: value  <= 0.56943088769912719727;
            RIGHT_4_4: value  <= 0.57886648178100585938;
            RIGHT_4_5: value  <= 0.55085647106170654297;
            RIGHT_4_6: value  <= 0.18572150170803070068;
            RIGHT_4_7: value  <= 0.21897700428962710295;
            RIGHT_4_8: value  <= 0.40438130497932428531;
            RIGHT_4_9: value  <= 0.54639732837677001953;
            RIGHT_4_10: value  <= 0.55909740924835205078;
            RIGHT_4_11: value  <= 0.26190540194511408023;
            RIGHT_4_12: value  <= 0.65352207422256469727;
            RIGHT_4_13: value  <= 0.55374461412429809570;
            RIGHT_4_14: value  <= 0.55447459220886230469;
            RIGHT_4_15: value  <= 0.30319759249687200375;
            RIGHT_4_16: value  <= 0.56465089321136474609;
            RIGHT_4_17: value  <= 0.54618209600448608398;
            RIGHT_4_18: value  <= 0.54592901468276977539;
            RIGHT_4_19: value  <= 0.28092199563980102539;
            RIGHT_4_20: value  <= 0.55038261413574218750;
            RIGHT_4_21: value  <= 0.33042821288108831235;
            RIGHT_4_22: value  <= 0.53789931535720825195;
            RIGHT_4_23: value  <= 0.22886039316654210873;
            RIGHT_4_24: value  <= 0.42529278993606567383;
            RIGHT_4_25: value  <= 0.53558301925659179688;
            RIGHT_4_26: value  <= 0.74425792694091796875;
            RIGHT_4_27: value  <= 0.25821250677108770200;
            RIGHT_4_28: value  <= 0.53610187768936157227;
            RIGHT_4_29: value  <= 0.45524680614471441098;
            RIGHT_4_30: value  <= 0.53440397977828979492;
            RIGHT_4_31: value  <= 0.56010431051254272461;
            RIGHT_4_32: value  <= 0.27688381075859069824;
            RIGHT_5_0: value  <= 0.61562412977218627930;
            RIGHT_5_1: value  <= 0.18323999643325811215;
            RIGHT_5_2: value  <= 0.57238161563873291016;
            RIGHT_5_3: value  <= 0.23772829771041870117;
            RIGHT_5_4: value  <= 0.58589351177215576172;
            RIGHT_5_5: value  <= 0.57941037416458129883;
            RIGHT_5_6: value  <= 0.24848650395870208740;
            RIGHT_5_7: value  <= 0.54842048883438110352;
            RIGHT_5_8: value  <= 0.60510927438735961914;
            RIGHT_5_9: value  <= 0.54412460327148437500;
            RIGHT_5_10: value  <= 0.23923380672931671143;
            RIGHT_5_11: value  <= 0.59646219015121459961;
            RIGHT_5_12: value  <= 0.15757469832897189055;
            RIGHT_5_13: value  <= 0.67484188079833984375;
            RIGHT_5_14: value  <= 0.54734510183334350586;
            RIGHT_5_15: value  <= 0.52271109819412231445;
            RIGHT_5_16: value  <= 0.61096358299255371094;
            RIGHT_5_17: value  <= 0.54040068387985229492;
            RIGHT_5_18: value  <= 0.22322730720043179597;
            RIGHT_5_19: value  <= 0.24536980688571929932;
            RIGHT_5_20: value  <= 0.53769302368164062500;
            RIGHT_5_21: value  <= 0.31556931138038640805;
            RIGHT_5_22: value  <= 0.65978652238845825195;
            RIGHT_5_23: value  <= 0.55052447319030761719;
            RIGHT_5_24: value  <= 0.18914650380611419678;
            RIGHT_5_25: value  <= 0.33442100882530212402;
            RIGHT_5_26: value  <= 0.23956120014190671053;
            RIGHT_5_27: value  <= 0.40222078561782842465;
            RIGHT_5_28: value  <= 0.45431908965110778809;
            RIGHT_5_29: value  <= 0.53577107191085815430;
            RIGHT_5_30: value  <= 0.71817511320114135742;
            RIGHT_5_31: value  <= 0.27917331457138061523;
            RIGHT_5_32: value  <= 0.39897239208221441098;
            RIGHT_5_33: value  <= 0.53006649017333984375;
            RIGHT_5_34: value  <= 0.52296727895736694336;
            RIGHT_5_35: value  <= 0.54534512758255004883;
            RIGHT_5_36: value  <= 0.44393768906593322754;
            RIGHT_5_37: value  <= 0.54893219470977783203;
            RIGHT_5_38: value  <= 0.42524749040603637695;
            RIGHT_5_39: value  <= 0.22926619648933410645;
            RIGHT_5_40: value  <= 0.40223899483680730649;
            RIGHT_5_41: value  <= 0.15361930429935460873;
            RIGHT_5_42: value  <= 0.52416062355041503906;
            RIGHT_5_43: value  <= 0.43251821398735051938;
            RIGHT_6_0: value  <= 0.14693309366703030672;
            RIGHT_6_1: value  <= 0.58964669704437255859;
            RIGHT_6_2: value  <= 0.17603619396686551180;
            RIGHT_6_3: value  <= 0.55960661172866821289;
            RIGHT_6_4: value  <= 0.57320362329483032227;
            RIGHT_6_5: value  <= 0.56230807304382324219;
            RIGHT_6_6: value  <= 0.56482332944869995117;
            RIGHT_6_7: value  <= 0.55046397447586059570;
            RIGHT_6_8: value  <= 0.57601428031921386719;
            RIGHT_6_9: value  <= 0.36597740650177001953;
            RIGHT_6_10: value  <= 0.59189391136169433594;
            RIGHT_6_11: value  <= 0.61831092834472656250;
            RIGHT_6_12: value  <= 0.31354010105133062192;
            RIGHT_6_13: value  <= 0.19166369736194610596;
            RIGHT_6_14: value  <= 0.66445910930633544922;
            RIGHT_6_15: value  <= 0.57093828916549682617;
            RIGHT_6_16: value  <= 0.56102699041366577148;
            RIGHT_6_17: value  <= 0.45803260803222661801;
            RIGHT_6_18: value  <= 0.29536840319633478336;
            RIGHT_6_19: value  <= 0.76190179586410522461;
            RIGHT_6_20: value  <= 0.17725290358066558838;
            RIGHT_6_21: value  <= 0.53407722711563110352;
            RIGHT_6_22: value  <= 0.60268038511276245117;
            RIGHT_6_23: value  <= 0.53243237733840942383;
            RIGHT_6_24: value  <= 0.53199452161788940430;
            RIGHT_6_25: value  <= 0.52103281021118164062;
            RIGHT_6_26: value  <= 0.34788420796394348145;
            RIGHT_6_27: value  <= 0.22576980292797088623;
            RIGHT_6_28: value  <= 0.52007079124450683594;
            RIGHT_6_29: value  <= 0.38201761245727539062;
            RIGHT_6_30: value  <= 0.66397482156753540039;
            RIGHT_6_31: value  <= 0.53823578357696533203;
            RIGHT_6_32: value  <= 0.42152971029281621762;
            RIGHT_6_33: value  <= 0.53863281011581420898;
            RIGHT_6_34: value  <= 0.68557357788085937500;
            RIGHT_6_35: value  <= 0.34674790501594537906;
            RIGHT_6_36: value  <= 0.43114539980888372250;
            RIGHT_6_37: value  <= 0.52249461412429809570;
            RIGHT_6_38: value  <= 0.54816448688507080078;
            RIGHT_6_39: value  <= 0.81826978921890258789;
            RIGHT_6_40: value  <= 0.52399927377700805664;
            RIGHT_6_41: value  <= 0.73781907558441162109;
            RIGHT_6_42: value  <= 0.44706439971923828125;
            RIGHT_6_43: value  <= 0.55379962921142578125;
            RIGHT_6_44: value  <= 0.53154432773590087891;
            RIGHT_6_45: value  <= 0.51387697458267211914;
            RIGHT_6_46: value  <= 0.33658531308174127750;
            RIGHT_6_47: value  <= 0.51626348495483398438;
            RIGHT_6_48: value  <= 0.44907060265541082211;
            RIGHT_6_49: value  <= 0.59855180978775024414;
            RIGHT_7_0: value  <= 0.66433167457580566406;
            RIGHT_7_1: value  <= 0.25185129046440130063;
            RIGHT_7_2: value  <= 0.23974630236625671387;
            RIGHT_7_3: value  <= 0.25291448831558227539;
            RIGHT_7_4: value  <= 0.55560797452926635742;
            RIGHT_7_5: value  <= 0.47628301382064819336;
            RIGHT_7_6: value  <= 0.28394040465354919434;
            RIGHT_7_7: value  <= 0.60063672065734863281;
            RIGHT_7_8: value  <= 0.27052891254425048828;
            RIGHT_7_9: value  <= 0.32622259855270391293;
            RIGHT_7_10: value  <= 0.41992568969726562500;
            RIGHT_7_11: value  <= 0.54348129034042358398;
            RIGHT_7_12: value  <= 0.23190039396286010742;
            RIGHT_7_13: value  <= 0.27082380652427667789;
            RIGHT_7_14: value  <= 0.58906257152557373047;
            RIGHT_7_15: value  <= 0.54199481010437011719;
            RIGHT_7_16: value  <= 0.27265900373458862305;
            RIGHT_7_17: value  <= 0.60172098875045776367;
            RIGHT_7_18: value  <= 0.14357580244541170988;
            RIGHT_7_19: value  <= 0.59299832582473754883;
            RIGHT_7_20: value  <= 0.30215978622436517886;
            RIGHT_7_21: value  <= 0.55320328474044799805;
            RIGHT_7_22: value  <= 0.33593991398811340332;
            RIGHT_7_23: value  <= 0.52304250001907348633;
            RIGHT_7_24: value  <= 0.10295289754867549548;
            RIGHT_7_25: value  <= 0.55582892894744873047;
            RIGHT_7_26: value  <= 0.18758599460124969482;
            RIGHT_7_27: value  <= 0.46796411275863647461;
            RIGHT_7_28: value  <= 0.43346709012985229492;
            RIGHT_7_29: value  <= 0.56502032279968261719;
            RIGHT_7_30: value  <= 0.52502560615539550781;
            RIGHT_7_31: value  <= 0.54459732770919799805;
            RIGHT_7_32: value  <= 0.62535631656646728516;
            RIGHT_7_33: value  <= 0.57000827789306640625;
            RIGHT_7_34: value  <= 0.65230387449264526367;
            RIGHT_7_35: value  <= 0.54281437397003173828;
            RIGHT_7_36: value  <= 0.39778938889503479004;
            RIGHT_7_37: value  <= 0.52195048332214355469;
            RIGHT_7_38: value  <= 0.55035740137100219727;
            RIGHT_7_39: value  <= 0.61223882436752319336;
            RIGHT_7_40: value  <= 0.51973849534988403320;
            RIGHT_7_41: value  <= 0.48931029438972467593;
            RIGHT_7_42: value  <= 0.54715752601623535156;
            RIGHT_7_43: value  <= 0.60739892721176147461;
            RIGHT_7_44: value  <= 0.46245330572128301450;
            RIGHT_7_45: value  <= 0.53066980838775634766;
            RIGHT_7_46: value  <= 0.25830659270286560059;
            RIGHT_7_47: value  <= 0.57354408502578735352;
            RIGHT_7_48: value  <= 0.44954448938369750977;
            RIGHT_7_49: value  <= 0.41381931304931640625;
            RIGHT_7_50: value  <= 0.43272399902343750000;
            RIGHT_8_0: value  <= 0.24822120368480679597;
            RIGHT_8_1: value  <= 0.23219659924507141113;
            RIGHT_8_2: value  <= 0.58149331808090209961;
            RIGHT_8_3: value  <= 0.58663117885589599609;
            RIGHT_8_4: value  <= 0.57913267612457275391;
            RIGHT_8_5: value  <= 0.56355422735214233398;
            RIGHT_8_6: value  <= 0.60547572374343872070;
            RIGHT_8_7: value  <= 0.27315109968185430356;
            RIGHT_8_8: value  <= 0.36385610699653631039;
            RIGHT_8_9: value  <= 0.54327291250228881836;
            RIGHT_8_10: value  <= 0.70698332786560058594;
            RIGHT_8_11: value  <= 0.52949970960617065430;
            RIGHT_8_12: value  <= 0.24977239966392519865;
            RIGHT_8_13: value  <= 0.57063561677932739258;
            RIGHT_8_14: value  <= 0.73947668075561523438;
            RIGHT_8_15: value  <= 0.24791529774665829744;
            RIGHT_8_16: value  <= 0.53389710187911987305;
            RIGHT_8_17: value  <= 0.53240692615509033203;
            RIGHT_8_18: value  <= 0.55345088243484497070;
            RIGHT_8_19: value  <= 0.65581941604614257812;
            RIGHT_8_20: value  <= 0.38102629780769348145;
            RIGHT_8_21: value  <= 0.57093858718872070312;
            RIGHT_8_22: value  <= 0.52595442533493041992;
            RIGHT_8_23: value  <= 0.57256120443344116211;
            RIGHT_8_24: value  <= 0.30444970726966857910;
            RIGHT_8_25: value  <= 0.55734348297119140625;
            RIGHT_8_26: value  <= 0.65188127756118774414;
            RIGHT_8_27: value  <= 0.55982369184494018555;
            RIGHT_8_28: value  <= 0.55618977546691894531;
            RIGHT_8_29: value  <= 0.53352999687194824219;
            RIGHT_8_30: value  <= 0.42213940620422357730;
            RIGHT_8_31: value  <= 0.21665850281715390291;
            RIGHT_8_32: value  <= 0.43546178936958307437;
            RIGHT_8_33: value  <= 0.35232171416282648257;
            RIGHT_8_34: value  <= 0.53384172916412353516;
            RIGHT_8_35: value  <= 0.37028178572654718570;
            RIGHT_8_36: value  <= 0.45836889743804931641;
            RIGHT_8_37: value  <= 0.39966610074043268375;
            RIGHT_8_38: value  <= 0.37774989008903497867;
            RIGHT_8_39: value  <= 0.51791828870773315430;
            RIGHT_8_40: value  <= 0.37001928687095642090;
            RIGHT_8_41: value  <= 0.56793761253356933594;
            RIGHT_8_42: value  <= 0.44809499382972717285;
            RIGHT_8_43: value  <= 0.53133869171142578125;
            RIGHT_8_44: value  <= 0.41293430328369140625;
            RIGHT_8_45: value  <= 0.56196212768554687500;
            RIGHT_8_46: value  <= 0.27205219864845281430;
            RIGHT_8_47: value  <= 0.66934937238693237305;
            RIGHT_8_48: value  <= 0.16372759640216830168;
            RIGHT_8_49: value  <= 0.29385319352149957828;
            RIGHT_8_50: value  <= 0.45322000980377197266;
            RIGHT_8_51: value  <= 0.35892319679260248355;
            RIGHT_8_52: value  <= 0.54411232471466064453;
            RIGHT_8_53: value  <= 0.40248918533325200864;
            RIGHT_8_54: value  <= 0.44226029515266418457;
            RIGHT_8_55: value  <= 0.17979049682617190276;
            RIGHT_9_0: value  <= 0.26265591382980352231;
            RIGHT_9_1: value  <= 0.57416272163391113281;
            RIGHT_9_2: value  <= 0.56266540288925170898;
            RIGHT_9_3: value  <= 0.19572949409484860506;
            RIGHT_9_4: value  <= 0.59925037622451782227;
            RIGHT_9_5: value  <= 0.60799038410186767578;
            RIGHT_9_6: value  <= 0.55769157409667968750;
            RIGHT_9_7: value  <= 0.55141717195510864258;
            RIGHT_9_8: value  <= 0.44770789146423339844;
            RIGHT_9_9: value  <= 0.26696211099624628238;
            RIGHT_9_10: value  <= 0.29888901114463811703;
            RIGHT_9_11: value  <= 0.51088631153106689453;
            RIGHT_9_12: value  <= 0.31203418970108032227;
            RIGHT_9_13: value  <= 0.56790757179260253906;
            RIGHT_9_14: value  <= 0.53448081016540527344;
            RIGHT_9_15: value  <= 0.53925681114196777344;
            RIGHT_9_16: value  <= 0.56927347183227539062;
            RIGHT_9_17: value  <= 0.54842978715896606445;
            RIGHT_9_18: value  <= 0.57560759782791137695;
            RIGHT_9_19: value  <= 0.47282311320304870605;
            RIGHT_9_20: value  <= 0.29323211312294011899;
            RIGHT_9_21: value  <= 0.42733490467071527652;
            RIGHT_9_22: value  <= 0.52064722776412963867;
            RIGHT_9_23: value  <= 0.16755220293998721037;
            RIGHT_9_24: value  <= 0.27776581048965448550;
            RIGHT_9_25: value  <= 0.48120489716529851743;
            RIGHT_9_26: value  <= 0.63491958379745483398;
            RIGHT_9_27: value  <= 0.53612488508224487305;
            RIGHT_9_28: value  <= 0.74096941947937011719;
            RIGHT_9_29: value  <= 0.54165017604827880859;
            RIGHT_9_30: value  <= 0.13117079436779019441;
            RIGHT_9_31: value  <= 0.25913399457931518555;
            RIGHT_9_32: value  <= 0.15823160111904138736;
            RIGHT_9_33: value  <= 0.43989789485931402035;
            RIGHT_9_34: value  <= 0.37080699205398559570;
            RIGHT_9_35: value  <= 0.55542111396789550781;
            RIGHT_9_36: value  <= 0.34111711382865911313;
            RIGHT_9_37: value  <= 0.43458628654479980469;
            RIGHT_9_38: value  <= 0.51937389373779296875;
            RIGHT_9_39: value  <= 0.47609439492225652524;
            RIGHT_9_40: value  <= 0.34113308787345891782;
            RIGHT_9_41: value  <= 0.55549472570419311523;
            RIGHT_9_42: value  <= 0.46974349021911621094;
            RIGHT_9_43: value  <= 0.39782929420471191406;
            RIGHT_9_44: value  <= 0.38455399870872497559;
            RIGHT_9_45: value  <= 0.53004968166351318359;
            RIGHT_9_46: value  <= 0.58288121223449707031;
            RIGHT_9_47: value  <= 0.52677577733993530273;
            RIGHT_9_48: value  <= 0.10236159712076189909;
            RIGHT_9_49: value  <= 0.43596929311752319336;
            RIGHT_9_50: value  <= 0.76060950756072998047;
            RIGHT_9_51: value  <= 0.18597120046615600586;
            RIGHT_9_52: value  <= 0.23320719599723818694;
            RIGHT_9_53: value  <= 0.32642349600791931152;
            RIGHT_9_54: value  <= 0.45332419872283941098;
            RIGHT_9_55: value  <= 0.54128098487854003906;
            RIGHT_9_56: value  <= 0.71386522054672241211;
            RIGHT_9_57: value  <= 0.54713201522827148438;
            RIGHT_9_58: value  <= 0.31304550170898437500;
            RIGHT_9_59: value  <= 0.34305301308631902524;
            RIGHT_9_60: value  <= 0.54686397314071655273;
            RIGHT_9_61: value  <= 0.53487008810043334961;
            RIGHT_9_62: value  <= 0.44926649332046508789;
            RIGHT_9_63: value  <= 0.52243089675903320312;
            RIGHT_9_64: value  <= 0.29933831095695501157;
            RIGHT_9_65: value  <= 0.44604998826980590820;
            RIGHT_9_66: value  <= 0.53881132602691650391;
            RIGHT_9_67: value  <= 0.48012199997901922055;
            RIGHT_9_68: value  <= 0.32614278793334960938;
            RIGHT_9_69: value  <= 0.57378298044204711914;
            RIGHT_9_70: value  <= 0.52338278293609619141;
            RIGHT_10_0: value  <= 0.68498080968856811523;
            RIGHT_10_1: value  <= 0.25378298759460449219;
            RIGHT_10_2: value  <= 0.28124240040779108218;
            RIGHT_10_3: value  <= 0.55442607402801513672;
            RIGHT_10_4: value  <= 0.54333502054214477539;
            RIGHT_10_5: value  <= 0.62207579612731933594;
            RIGHT_10_6: value  <= 0.29923579096794128418;
            RIGHT_10_7: value  <= 0.54116767644882202148;
            RIGHT_10_8: value  <= 0.53645849227905273438;
            RIGHT_10_9: value  <= 0.57296061515808105469;
            RIGHT_10_10: value  <= 0.52582687139511108398;
            RIGHT_10_11: value  <= 0.38511589169502258301;
            RIGHT_10_12: value  <= 0.36365869641304021664;
            RIGHT_10_13: value  <= 0.53775602579116821289;
            RIGHT_10_14: value  <= 0.55724847316741943359;
            RIGHT_10_15: value  <= 0.45325040817260742188;
            RIGHT_10_16: value  <= 0.29325398802757257632;
            RIGHT_10_17: value  <= 0.53300672769546508789;
            RIGHT_10_18: value  <= 0.51193618774414062500;
            RIGHT_10_19: value  <= 0.70083981752395629883;
            RIGHT_10_20: value  <= 0.51041620969772338867;
            RIGHT_10_21: value  <= 0.13061730563640588931;
            RIGHT_10_22: value  <= 0.54398590326309204102;
            RIGHT_10_23: value  <= 0.76875698566436767578;
            RIGHT_10_24: value  <= 0.32409390807151788882;
            RIGHT_10_25: value  <= 0.52304041385650634766;
            RIGHT_10_26: value  <= 0.55179458856582641602;
            RIGHT_10_27: value  <= 0.61317539215087890625;
            RIGHT_10_28: value  <= 0.52807378768920898438;
            RIGHT_10_29: value  <= 0.48560309410095220395;
            RIGHT_10_30: value  <= 0.52560812234878540039;
            RIGHT_10_31: value  <= 0.62772971391677856445;
            RIGHT_10_32: value  <= 0.45750290155410772153;
            RIGHT_10_33: value  <= 0.54694122076034545898;
            RIGHT_10_34: value  <= 0.67687010765075683594;
            RIGHT_10_35: value  <= 0.37917000055313110352;
            RIGHT_10_36: value  <= 0.58734762668609619141;
            RIGHT_10_37: value  <= 0.55852657556533813477;
            RIGHT_10_38: value  <= 0.46035489439964288882;
            RIGHT_10_39: value  <= 0.59002387523651123047;
            RIGHT_10_40: value  <= 0.18088449537754058838;
            RIGHT_10_41: value  <= 0.37178671360015869141;
            RIGHT_10_42: value  <= 0.51488637924194335938;
            RIGHT_10_43: value  <= 0.47387400269508361816;
            RIGHT_10_44: value  <= 0.63031142950057983398;
            RIGHT_10_45: value  <= 0.37021011114120477847;
            RIGHT_10_46: value  <= 0.51014107465744018555;
            RIGHT_10_47: value  <= 0.51687937974929809570;
            RIGHT_10_48: value  <= 0.63138538599014282227;
            RIGHT_10_49: value  <= 0.53773492574691772461;
            RIGHT_10_50: value  <= 0.36642369627952581235;
            RIGHT_10_51: value  <= 0.35415500402450561523;
            RIGHT_10_52: value  <= 0.56672430038452148438;
            RIGHT_10_53: value  <= 0.51986688375473022461;
            RIGHT_10_54: value  <= 0.50281071662902832031;
            RIGHT_10_55: value  <= 0.62227207422256469727;
            RIGHT_10_56: value  <= 0.51378047466278076172;
            RIGHT_10_57: value  <= 0.37217769026756292172;
            RIGHT_10_58: value  <= 0.46852919459342962094;
            RIGHT_10_59: value  <= 0.42403739690780639648;
            RIGHT_10_60: value  <= 0.35013249516487121582;
            RIGHT_10_61: value  <= 0.47265690565109247379;
            RIGHT_10_62: value  <= 0.07574920356273649735;
            RIGHT_10_63: value  <= 0.55385738611221313477;
            RIGHT_10_64: value  <= 0.53596121072769165039;
            RIGHT_10_65: value  <= 0.46493428945541381836;
            RIGHT_10_66: value  <= 0.43471878767013549805;
            RIGHT_10_67: value  <= 0.23155799508094790373;
            RIGHT_10_68: value  <= 0.29773768782615661621;
            RIGHT_10_69: value  <= 0.48615050315856928043;
            RIGHT_10_70: value  <= 0.52298247814178466797;
            RIGHT_10_71: value  <= 0.52101737260818481445;
            RIGHT_10_72: value  <= 0.65850979089736938477;
            RIGHT_10_73: value  <= 0.51989167928695678711;
            RIGHT_10_74: value  <= 0.46513590216636657715;
            RIGHT_10_75: value  <= 0.58985459804534912109;
            RIGHT_10_76: value  <= 0.53660178184509277344;
            RIGHT_10_77: value  <= 0.83152848482131958008;
            RIGHT_10_78: value  <= 0.53705602884292602539;
            RIGHT_10_79: value  <= 0.59673351049423217773;
            RIGHT_11_0: value  <= 0.30545330047607421875;
            RIGHT_11_1: value  <= 0.31555780768394470215;
            RIGHT_11_2: value  <= 0.56929117441177368164;
            RIGHT_11_3: value  <= 0.59349310398101806641;
            RIGHT_11_4: value  <= 0.54747921228408813477;
            RIGHT_11_5: value  <= 0.56675457954406738281;
            RIGHT_11_6: value  <= 0.58454728126525878906;
            RIGHT_11_7: value  <= 0.55228072404861450195;
            RIGHT_11_8: value  <= 0.53754240274429321289;
            RIGHT_11_9: value  <= 0.54989522695541381836;
            RIGHT_11_10: value  <= 0.63137108087539672852;
            RIGHT_11_11: value  <= 0.40526661276817321777;
            RIGHT_11_12: value  <= 0.23186540603637700864;
            RIGHT_11_13: value  <= 0.52415257692337036133;
            RIGHT_11_14: value  <= 0.36771959066390991211;
            RIGHT_11_15: value  <= 0.55424308776855468750;
            RIGHT_11_16: value  <= 0.53009599447250366211;
            RIGHT_11_17: value  <= 0.57954281568527221680;
            RIGHT_11_18: value  <= 0.52920591831207275391;
            RIGHT_11_19: value  <= 0.47481718659400939941;
            RIGHT_11_20: value  <= 0.55768972635269165039;
            RIGHT_11_21: value  <= 0.52867668867111206055;
            RIGHT_11_22: value  <= 0.34862980246543878726;
            RIGHT_11_23: value  <= 0.46768361330032348633;
            RIGHT_11_24: value  <= 0.46607351303100591489;
            RIGHT_11_25: value  <= 0.53512877225875854492;
            RIGHT_11_26: value  <= 0.32896101474761957340;
            RIGHT_11_27: value  <= 0.47543001174926757812;
            RIGHT_11_28: value  <= 0.53605020046234130859;
            RIGHT_11_29: value  <= 0.35520640015602111816;
            RIGHT_11_30: value  <= 0.12564620375633239746;
            RIGHT_11_31: value  <= 0.16258180141448980160;
            RIGHT_11_32: value  <= 0.45841971039772028140;
            RIGHT_11_33: value  <= 0.34946969151496892758;
            RIGHT_11_34: value  <= 0.51602262258529663086;
            RIGHT_11_35: value  <= 0.57679080963134765625;
            RIGHT_11_36: value  <= 0.53477007150650024414;
            RIGHT_11_37: value  <= 0.63872468471527099609;
            RIGHT_11_38: value  <= 0.41203960776329040527;
            RIGHT_11_39: value  <= 0.70898222923278808594;
            RIGHT_11_40: value  <= 0.28952449560165410825;
            RIGHT_11_41: value  <= 0.52196067571640014648;
            RIGHT_11_42: value  <= 0.49998161196708679199;
            RIGHT_11_43: value  <= 0.40296629071235662289;
            RIGHT_11_44: value  <= 0.58662968873977661133;
            RIGHT_11_45: value  <= 0.49190279841423040219;
            RIGHT_11_46: value  <= 0.53487390279769897461;
            RIGHT_11_47: value  <= 0.61299049854278564453;
            RIGHT_11_48: value  <= 0.34234538674354547672;
            RIGHT_11_49: value  <= 0.58243042230606079102;
            RIGHT_11_50: value  <= 0.28561499714851379395;
            RIGHT_11_51: value  <= 0.59585297107696533203;
            RIGHT_11_52: value  <= 0.47414121031761169434;
            RIGHT_11_53: value  <= 0.53372788429260253906;
            RIGHT_11_54: value  <= 0.67258632183074951172;
            RIGHT_11_55: value  <= 0.28456708788871770688;
            RIGHT_11_56: value  <= 0.57185977697372436523;
            RIGHT_11_57: value  <= 0.28048470616340642758;
            RIGHT_11_58: value  <= 0.33145239949226379395;
            RIGHT_11_59: value  <= 0.62769711017608642578;
            RIGHT_11_60: value  <= 0.20171439647674560547;
            RIGHT_11_61: value  <= 0.48766410350799560547;
            RIGHT_11_62: value  <= 0.58812642097473144531;
            RIGHT_11_63: value  <= 0.52860087156295776367;
            RIGHT_11_64: value  <= 0.45880940556526178531;
            RIGHT_11_65: value  <= 0.54859781265258789062;
            RIGHT_11_66: value  <= 0.52541971206665039062;
            RIGHT_11_67: value  <= 0.54540151357650756836;
            RIGHT_11_68: value  <= 0.44858568906784057617;
            RIGHT_11_69: value  <= 0.39253529906272888184;
            RIGHT_11_70: value  <= 0.45885840058326721191;
            RIGHT_11_71: value  <= 0.53698569536209106445;
            RIGHT_11_72: value  <= 0.37057501077651977539;
            RIGHT_11_73: value  <= 0.64527308940887451172;
            RIGHT_11_74: value  <= 0.40646770596504211426;
            RIGHT_11_75: value  <= 0.52947628498077392578;
            RIGHT_11_76: value  <= 0.51449728012084960938;
            RIGHT_11_77: value  <= 0.48520979285240167789;
            RIGHT_11_78: value  <= 0.41530540585517877750;
            RIGHT_11_79: value  <= 0.45663040876388549805;
            RIGHT_11_80: value  <= 0.51881599426269531250;
            RIGHT_11_81: value  <= 0.22026319801807400789;
            RIGHT_11_82: value  <= 0.50603431463241577148;
            RIGHT_11_83: value  <= 0.11850229650735860654;
            RIGHT_11_84: value  <= 0.68261492252349853516;
            RIGHT_11_85: value  <= 0.52250087261199951172;
            RIGHT_11_86: value  <= 0.50808018445968627930;
            RIGHT_11_87: value  <= 0.47904640436172490903;
            RIGHT_11_88: value  <= 0.15635989606380459871;
            RIGHT_11_89: value  <= 0.72305107116699218750;
            RIGHT_11_90: value  <= 0.50987982749938964844;
            RIGHT_11_91: value  <= 0.67709028720855712891;
            RIGHT_11_92: value  <= 0.50810241699218750000;
            RIGHT_11_93: value  <= 0.48103410005569458008;
            RIGHT_11_94: value  <= 0.52354729175567626953;
            RIGHT_11_95: value  <= 0.49192130565643310547;
            RIGHT_11_96: value  <= 0.60821849107742309570;
            RIGHT_11_97: value  <= 0.32924321293830871582;
            RIGHT_11_98: value  <= 0.45949959754943847656;
            RIGHT_11_99: value  <= 0.57672828435897827148;
            RIGHT_11_100: value  <= 0.26350161433219909668;
            RIGHT_11_101: value  <= 0.52789801359176635742;
            RIGHT_11_102: value  <= 0.55175000429153442383;
            RIGHT_12_0: value  <= 0.63352262973785400391;
            RIGHT_12_1: value  <= 0.34774878621101379395;
            RIGHT_12_2: value  <= 0.55821180343627929688;
            RIGHT_12_3: value  <= 0.59300708770751953125;
            RIGHT_12_4: value  <= 0.33479958772659301758;
            RIGHT_12_5: value  <= 0.55086308717727661133;
            RIGHT_12_6: value  <= 0.36990478634834289551;
            RIGHT_12_7: value  <= 0.54379111528396606445;
            RIGHT_12_8: value  <= 0.17957249283790591154;
            RIGHT_12_9: value  <= 0.44468268752098077945;
            RIGHT_12_10: value  <= 0.53469717502593994141;
            RIGHT_12_11: value  <= 0.53311979770660400391;
            RIGHT_12_12: value  <= 0.45880630612373352051;
            RIGHT_12_13: value  <= 0.22744719684123990144;
            RIGHT_12_14: value  <= 0.38150069117546081543;
            RIGHT_12_15: value  <= 0.25437268614768981934;
            RIGHT_12_16: value  <= 0.34063041210174560547;
            RIGHT_12_17: value  <= 0.54205721616744995117;
            RIGHT_12_18: value  <= 0.56601101160049438477;
            RIGHT_12_19: value  <= 0.39406880736351007632;
            RIGHT_12_20: value  <= 0.71185618638992309570;
            RIGHT_12_21: value  <= 0.53221440315246582031;
            RIGHT_12_22: value  <= 0.51220291852951049805;
            RIGHT_12_23: value  <= 0.64554882049560546875;
            RIGHT_12_24: value  <= 0.23616339266300198640;
            RIGHT_12_25: value  <= 0.44766610860824590512;
            RIGHT_12_26: value  <= 0.51022082567214965820;
            RIGHT_12_27: value  <= 0.15359309315681460295;
            RIGHT_12_28: value  <= 0.36246618628501892090;
            RIGHT_12_29: value  <= 0.48455920815467828922;
            RIGHT_12_30: value  <= 0.58241981267929077148;
            RIGHT_12_31: value  <= 0.14394679665565490723;
            RIGHT_12_32: value  <= 0.52870452404022216797;
            RIGHT_12_33: value  <= 0.61220401525497436523;
            RIGHT_12_34: value  <= 0.50455862283706665039;
            RIGHT_12_35: value  <= 0.47947341203689580746;
            RIGHT_12_36: value  <= 0.24985109269618990813;
            RIGHT_12_37: value  <= 0.37095320224761957340;
            RIGHT_12_38: value  <= 0.50816917419433593750;
            RIGHT_12_39: value  <= 0.47836089134216308594;
            RIGHT_12_40: value  <= 0.44998261332511901855;
            RIGHT_12_41: value  <= 0.54193347692489624023;
            RIGHT_12_42: value  <= 0.12157420068979260530;
            RIGHT_12_43: value  <= 0.53818839788436889648;
            RIGHT_12_44: value  <= 0.57034862041473388672;
            RIGHT_12_45: value  <= 0.55475491285324096680;
            RIGHT_12_46: value  <= 0.50970828533172607422;
            RIGHT_12_47: value  <= 0.43030360341072082520;
            RIGHT_12_48: value  <= 0.69820040464401245117;
            RIGHT_12_49: value  <= 0.22690680623054498843;
            RIGHT_12_50: value  <= 0.45379561185836791992;
            RIGHT_12_51: value  <= 0.27404838800430297852;
            RIGHT_12_52: value  <= 0.50717329978942871094;
            RIGHT_12_53: value  <= 0.61198681592941284180;
            RIGHT_12_54: value  <= 0.20282049477100369539;
            RIGHT_12_55: value  <= 0.54308217763900756836;
            RIGHT_12_56: value  <= 0.67793232202529907227;
            RIGHT_12_57: value  <= 0.34314650297164922543;
            RIGHT_12_58: value  <= 0.50032228231430053711;
            RIGHT_12_59: value  <= 0.15906329452991491147;
            RIGHT_12_60: value  <= 0.46480441093444818668;
            RIGHT_12_61: value  <= 0.39231911301612848453;
            RIGHT_12_62: value  <= 0.46291279792785650082;
            RIGHT_12_63: value  <= 0.52061259746551513672;
            RIGHT_12_64: value  <= 0.30538770556449890137;
            RIGHT_12_65: value  <= 0.51690948009490966797;
            RIGHT_12_66: value  <= 0.42308250069618230649;
            RIGHT_12_67: value  <= 0.40797919034957891293;
            RIGHT_12_68: value  <= 0.45744091272354131528;
            RIGHT_12_69: value  <= 0.51950198411941528320;
            RIGHT_12_70: value  <= 0.50434887409210205078;
            RIGHT_12_71: value  <= 0.47575059533119201660;
            RIGHT_12_72: value  <= 0.50650137662887573242;
            RIGHT_12_73: value  <= 0.56658387184143066406;
            RIGHT_12_74: value  <= 0.55868571996688842773;
            RIGHT_12_75: value  <= 0.48127061128616327457;
            RIGHT_12_76: value  <= 0.52870899438858032227;
            RIGHT_12_77: value  <= 0.59240859746932983398;
            RIGHT_12_78: value  <= 0.06915248185396190295;
            RIGHT_12_79: value  <= 0.49340128898620611020;
            RIGHT_12_80: value  <= 0.58934777975082397461;
            RIGHT_12_81: value  <= 0.53962701559066772461;
            RIGHT_12_82: value  <= 0.50683307647705078125;
            RIGHT_12_83: value  <= 0.42435330152511602231;
            RIGHT_12_84: value  <= 0.45400860905647277832;
            RIGHT_12_85: value  <= 0.30261999368667602539;
            RIGHT_12_86: value  <= 0.25576829910278320312;
            RIGHT_12_87: value  <= 0.58618277311325073242;
            RIGHT_12_88: value  <= 0.15271779894828799162;
            RIGHT_12_89: value  <= 0.48906040191650390625;
            RIGHT_12_90: value  <= 0.45146000385284418277;
            RIGHT_12_91: value  <= 0.54009538888931274414;
            RIGHT_12_92: value  <= 0.50740778446197509766;
            RIGHT_12_93: value  <= 0.54025697708129882812;
            RIGHT_12_94: value  <= 0.45950970053672790527;
            RIGHT_12_95: value  <= 0.45005279779434198550;
            RIGHT_12_96: value  <= 0.53107571601867675781;
            RIGHT_12_97: value  <= 0.47561758756637567691;
            RIGHT_12_98: value  <= 0.54510641098022460938;
            RIGHT_12_99: value  <= 0.48247399926185607910;
            RIGHT_12_100: value  <= 0.51573359966278076172;
            RIGHT_12_101: value  <= 0.71599560976028442383;
            RIGHT_12_102: value  <= 0.46192750334739690610;
            RIGHT_12_103: value  <= 0.24506139755249020662;
            RIGHT_12_104: value  <= 0.63940370082855224609;
            RIGHT_12_105: value  <= 0.54836612939834594727;
            RIGHT_12_106: value  <= 0.27014800906181341000;
            RIGHT_12_107: value  <= 0.53874611854553222656;
            RIGHT_12_108: value  <= 0.37194138765335077457;
            RIGHT_12_109: value  <= 0.68951261043548583984;
            RIGHT_12_110: value  <= 0.39180809259414667300;
            RIGHT_13_0: value  <= 0.71425348520278930664;
            RIGHT_13_1: value  <= 0.60900169610977172852;
            RIGHT_13_2: value  <= 0.59879022836685180664;
            RIGHT_13_3: value  <= 0.56972408294677734375;
            RIGHT_13_4: value  <= 0.55316567420959472656;
            RIGHT_13_5: value  <= 0.56726312637329101562;
            RIGHT_13_6: value  <= 0.53887271881103515625;
            RIGHT_13_7: value  <= 0.54987788200378417969;
            RIGHT_13_8: value  <= 0.27628791332244867496;
            RIGHT_13_9: value  <= 0.52592468261718750000;
            RIGHT_13_10: value  <= 0.40736979246139531918;
            RIGHT_13_11: value  <= 0.54158622026443481445;
            RIGHT_13_12: value  <= 0.35031560063362121582;
            RIGHT_13_13: value  <= 0.34111958742141718082;
            RIGHT_13_14: value  <= 0.53353762626647949219;
            RIGHT_13_15: value  <= 0.55365538597106933594;
            RIGHT_13_16: value  <= 0.52480888366699218750;
            RIGHT_13_17: value  <= 0.66060417890548706055;
            RIGHT_13_18: value  <= 0.52876251935958862305;
            RIGHT_13_19: value  <= 0.47499281167984008789;
            RIGHT_13_20: value  <= 0.50989967584609985352;
            RIGHT_13_21: value  <= 0.58811670541763305664;
            RIGHT_13_22: value  <= 0.90897941589355468750;
            RIGHT_13_23: value  <= 0.55778372287750244141;
            RIGHT_13_24: value  <= 0.65808779001235961914;
            RIGHT_13_25: value  <= 0.39758789539337158203;
            RIGHT_13_26: value  <= 0.36054858565330510922;
            RIGHT_13_27: value  <= 0.17967459559440610017;
            RIGHT_13_28: value  <= 0.51140302419662475586;
            RIGHT_13_29: value  <= 0.66082191467285156250;
            RIGHT_13_30: value  <= 0.44368579983711242676;
            RIGHT_13_31: value  <= 0.40540221333503717593;
            RIGHT_13_32: value  <= 0.32734549045562738590;
            RIGHT_13_33: value  <= 0.49757811427116388492;
            RIGHT_13_34: value  <= 0.35609039664268488101;
            RIGHT_13_35: value  <= 0.58164817094802856445;
            RIGHT_13_36: value  <= 0.34464201331138610840;
            RIGHT_13_37: value  <= 0.74721592664718627930;
            RIGHT_13_38: value  <= 0.64017212390899658203;
            RIGHT_13_39: value  <= 0.35552209615707397461;
            RIGHT_13_40: value  <= 0.57727241516113281250;
            RIGHT_13_41: value  <= 0.52929002046585083008;
            RIGHT_13_42: value  <= 0.16755819320678710938;
            RIGHT_13_43: value  <= 0.70856010913848876953;
            RIGHT_13_44: value  <= 0.21624700725078579988;
            RIGHT_13_45: value  <= 0.52513718605041503906;
            RIGHT_13_46: value  <= 0.41978681087493902035;
            RIGHT_13_47: value  <= 0.54296958446502685547;
            RIGHT_13_48: value  <= 0.25145179033279418945;
            RIGHT_13_49: value  <= 0.48496189713478088379;
            RIGHT_13_50: value  <= 0.53944462537765502930;
            RIGHT_13_51: value  <= 0.45691820979118352719;
            RIGHT_13_52: value  <= 0.28022980690002441406;
            RIGHT_13_53: value  <= 0.46361210942268371582;
            RIGHT_13_54: value  <= 0.52546602487564086914;
            RIGHT_13_55: value  <= 0.40820831060409551450;
            RIGHT_13_56: value  <= 0.58065170049667358398;
            RIGHT_13_57: value  <= 0.51827752590179443359;
            RIGHT_13_58: value  <= 0.34561741352081298828;
            RIGHT_13_59: value  <= 0.59424138069152832031;
            RIGHT_13_60: value  <= 0.70248460769653320312;
            RIGHT_13_61: value  <= 0.37689670920372009277;
            RIGHT_13_62: value  <= 0.54574978351593017578;
            RIGHT_13_63: value  <= 0.51549088954925537109;
            RIGHT_13_64: value  <= 0.27918958663940429688;
            RIGHT_13_65: value  <= 0.47563329339027410336;
            RIGHT_13_66: value  <= 0.40926858782768249512;
            RIGHT_13_67: value  <= 0.52855509519577026367;
            RIGHT_13_68: value  <= 0.46528089046478271484;
            RIGHT_13_69: value  <= 0.45027598738670349121;
            RIGHT_13_70: value  <= 0.45725551247596740723;
            RIGHT_13_71: value  <= 0.51816147565841674805;
            RIGHT_13_72: value  <= 0.51949840784072875977;
            RIGHT_13_73: value  <= 0.48518198728561401367;
            RIGHT_13_74: value  <= 0.55198061466217041016;
            RIGHT_13_75: value  <= 0.42085149884223937988;
            RIGHT_13_76: value  <= 0.45606550574302667789;
            RIGHT_13_77: value  <= 0.22582270205020910092;
            RIGHT_13_78: value  <= 0.51567047834396362305;
            RIGHT_13_79: value  <= 0.66899412870407104492;
            RIGHT_13_80: value  <= 0.52510780096054077148;
            RIGHT_13_81: value  <= 0.49663299322128301450;
            RIGHT_13_82: value  <= 0.50611138343811035156;
            RIGHT_13_83: value  <= 0.42380660772323608398;
            RIGHT_13_84: value  <= 0.54977869987487792969;
            RIGHT_13_85: value  <= 0.56642740964889526367;
            RIGHT_13_86: value  <= 0.44631358981132507324;
            RIGHT_13_87: value  <= 0.52210032939910888672;
            RIGHT_13_88: value  <= 0.50063651800155639648;
            RIGHT_13_89: value  <= 0.12822559475898739900;
            RIGHT_13_90: value  <= 0.73639607429504394531;
            RIGHT_13_91: value  <= 0.55189967155456542969;
            RIGHT_13_92: value  <= 0.36851361393928527832;
            RIGHT_13_93: value  <= 0.47162809967994689941;
            RIGHT_13_94: value  <= 0.37761849164962768555;
            RIGHT_13_95: value  <= 0.51983469724655151367;
            RIGHT_13_96: value  <= 0.38389080762863159180;
            RIGHT_13_97: value  <= 0.57552242279052734375;
            RIGHT_13_98: value  <= 0.51667708158493041992;
            RIGHT_13_99: value  <= 0.64597177505493164062;
            RIGHT_13_100: value  <= 0.60102558135986328125;
            RIGHT_13_101: value  <= 0.54932558536529541016;
            RIGHT_14_0: value  <= 0.37438011169433588199;
            RIGHT_14_1: value  <= 0.34377971291542047672;
            RIGHT_14_2: value  <= 0.59082162380218505859;
            RIGHT_14_3: value  <= 0.28735581040382390805;
            RIGHT_14_4: value  <= 0.54310190677642822266;
            RIGHT_14_5: value  <= 0.57413887977600097656;
            RIGHT_14_6: value  <= 0.34628450870513921567;
            RIGHT_14_7: value  <= 0.54295092821121215820;
            RIGHT_14_8: value  <= 0.53518110513687133789;
            RIGHT_14_9: value  <= 0.57002341747283935547;
            RIGHT_14_10: value  <= 0.33668708801269531250;
            RIGHT_14_11: value  <= 0.62573361396789550781;
            RIGHT_14_12: value  <= 0.51294529438018798828;
            RIGHT_14_13: value  <= 0.41550621390342712402;
            RIGHT_14_14: value  <= 0.58045381307601928711;
            RIGHT_14_15: value  <= 0.52026861906051635742;
            RIGHT_14_16: value  <= 0.35856771469116210938;
            RIGHT_14_17: value  <= 0.59415858983993530273;
            RIGHT_14_18: value  <= 0.50887960195541381836;
            RIGHT_14_19: value  <= 0.68410611152648925781;
            RIGHT_14_20: value  <= 0.37484970688819890805;
            RIGHT_14_21: value  <= 0.38538050651550287418;
            RIGHT_14_22: value  <= 0.53409588336944580078;
            RIGHT_14_23: value  <= 0.60599899291992187500;
            RIGHT_14_24: value  <= 0.60124689340591430664;
            RIGHT_14_25: value  <= 0.18403880298137670346;
            RIGHT_14_26: value  <= 0.44098970293998718262;
            RIGHT_14_27: value  <= 0.55892372131347656250;
            RIGHT_14_28: value  <= 0.20626190304756170102;
            RIGHT_14_29: value  <= 0.41926109790802001953;
            RIGHT_14_30: value  <= 0.40033689141273498535;
            RIGHT_14_31: value  <= 0.54441910982131958008;
            RIGHT_14_32: value  <= 0.39449059963226318359;
            RIGHT_14_33: value  <= 0.41927140951156621762;
            RIGHT_14_34: value  <= 0.46049609780311578922;
            RIGHT_14_35: value  <= 0.29268300533294677734;
            RIGHT_14_36: value  <= 0.73074632883071899414;
            RIGHT_14_37: value  <= 0.54150652885437011719;
            RIGHT_14_38: value  <= 0.56040412187576293945;
            RIGHT_14_39: value  <= 0.52931827306747436523;
            RIGHT_14_40: value  <= 0.46218210458755487613;
            RIGHT_14_41: value  <= 0.54204392433166503906;
            RIGHT_14_42: value  <= 0.50378918647766113281;
            RIGHT_14_43: value  <= 0.56139731407165527344;
            RIGHT_14_44: value  <= 0.59261232614517211914;
            RIGHT_14_45: value  <= 0.37283858656883239746;
            RIGHT_14_46: value  <= 0.29756438732147222348;
            RIGHT_14_47: value  <= 0.48245379328727722168;
            RIGHT_14_48: value  <= 0.64147979021072387695;
            RIGHT_14_49: value  <= 0.34299948811531072446;
            RIGHT_14_50: value  <= 0.50133150815963745117;
            RIGHT_14_51: value  <= 0.46974050998687738590;
            RIGHT_14_52: value  <= 0.64365047216415405273;
            RIGHT_14_53: value  <= 0.60438942909240722656;
            RIGHT_14_54: value  <= 0.32318168878555297852;
            RIGHT_14_55: value  <= 0.52009809017181396484;
            RIGHT_14_56: value  <= 0.38156008720397949219;
            RIGHT_14_57: value  <= 0.46889019012451171875;
            RIGHT_14_58: value  <= 0.62874001264572143555;
            RIGHT_14_59: value  <= 0.33036559820175170898;
            RIGHT_14_60: value  <= 0.50054347515106201172;
            RIGHT_14_61: value  <= 0.43251338601112371274;
            RIGHT_14_62: value  <= 0.54477912187576293945;
            RIGHT_14_63: value  <= 0.67786490917205810547;
            RIGHT_14_64: value  <= 0.36121138930320739746;
            RIGHT_14_65: value  <= 0.32502880692482000180;
            RIGHT_14_66: value  <= 0.66659259796142578125;
            RIGHT_14_67: value  <= 0.38836041092872619629;
            RIGHT_14_68: value  <= 0.73018449544906616211;
            RIGHT_14_69: value  <= 0.54649841785430908203;
            RIGHT_14_70: value  <= 0.50895309448242187500;
            RIGHT_14_71: value  <= 0.49407958984375000000;
            RIGHT_14_72: value  <= 0.78787708282470703125;
            RIGHT_14_73: value  <= 0.27484980225563049316;
            RIGHT_14_74: value  <= 0.40419089794158941098;
            RIGHT_14_75: value  <= 0.48152831196784967593;
            RIGHT_14_76: value  <= 0.70289808511734008789;
            RIGHT_14_77: value  <= 0.53046840429306030273;
            RIGHT_14_78: value  <= 0.46888920664787292480;
            RIGHT_14_79: value  <= 0.55734640359878540039;
            RIGHT_14_80: value  <= 0.52639877796173095703;
            RIGHT_14_81: value  <= 0.53872710466384887695;
            RIGHT_14_82: value  <= 0.74472510814666748047;
            RIGHT_14_83: value  <= 0.55919218063354492188;
            RIGHT_14_84: value  <= 0.46769270300865167789;
            RIGHT_14_85: value  <= 0.33081620931625371762;
            RIGHT_14_86: value  <= 0.33090591430664062500;
            RIGHT_14_87: value  <= 0.60783427953720092773;
            RIGHT_14_88: value  <= 0.58639198541641235352;
            RIGHT_14_89: value  <= 0.42085230350494390317;
            RIGHT_14_90: value  <= 0.40006220340728759766;
            RIGHT_14_91: value  <= 0.42596429586410522461;
            RIGHT_14_92: value  <= 0.33508691191673278809;
            RIGHT_14_93: value  <= 0.71473097801208496094;
            RIGHT_14_94: value  <= 0.50837898254394531250;
            RIGHT_14_95: value  <= 0.50217670202255249023;
            RIGHT_14_96: value  <= 0.55225551128387451172;
            RIGHT_14_97: value  <= 0.53900748491287231445;
            RIGHT_14_98: value  <= 0.75043660402297973633;
            RIGHT_14_99: value  <= 0.55383628606796264648;
            RIGHT_14_100: value  <= 0.45297130942344671078;
            RIGHT_14_101: value  <= 0.54733997583389282227;
            RIGHT_14_102: value  <= 0.57979941368103027344;
            RIGHT_14_103: value  <= 0.44324448704719537906;
            RIGHT_14_104: value  <= 0.63642418384552001953;
            RIGHT_14_105: value  <= 0.59144157171249389648;
            RIGHT_14_106: value  <= 0.38859179615974431821;
            RIGHT_14_107: value  <= 0.37449419498443597965;
            RIGHT_14_108: value  <= 0.56146162748336791992;
            RIGHT_14_109: value  <= 0.51855427026748657227;
            RIGHT_14_110: value  <= 0.56828498840332031250;
            RIGHT_14_111: value  <= 0.23793940246105191316;
            RIGHT_14_112: value  <= 0.44664269685745239258;
            RIGHT_14_113: value  <= 0.52510571479797363281;
            RIGHT_14_114: value  <= 0.33975180983543401547;
            RIGHT_14_115: value  <= 0.48459240794181818179;
            RIGHT_14_116: value  <= 0.34541139006614690610;
            RIGHT_14_117: value  <= 0.51886677742004394531;
            RIGHT_14_118: value  <= 0.56557738780975341797;
            RIGHT_14_119: value  <= 0.49592170119285577945;
            RIGHT_14_120: value  <= 0.50322318077087402344;
            RIGHT_14_121: value  <= 0.27551281452178960629;
            RIGHT_14_122: value  <= 0.52145522832870483398;
            RIGHT_14_123: value  <= 0.45111650228500371762;
            RIGHT_14_124: value  <= 0.73315447568893432617;
            RIGHT_14_125: value  <= 0.41015630960464477539;
            RIGHT_14_126: value  <= 0.12729619443416601010;
            RIGHT_14_127: value  <= 0.51656562089920043945;
            RIGHT_14_128: value  <= 0.46842318773269647769;
            RIGHT_14_129: value  <= 0.47889319062232971191;
            RIGHT_14_130: value  <= 0.52205038070678710938;
            RIGHT_14_131: value  <= 0.52396631240844726562;
            RIGHT_14_132: value  <= 0.24252149462699890137;
            RIGHT_14_133: value  <= 0.47585740685462951660;
            RIGHT_14_134: value  <= 0.52635979652404785156;
            RIGHT_15_0: value  <= 0.62405228614807128906;
            RIGHT_15_1: value  <= 0.69429391622543334961;
            RIGHT_15_2: value  <= 0.59007328748703002930;
            RIGHT_15_3: value  <= 0.53005450963973999023;
            RIGHT_15_4: value  <= 0.31031790375709528140;
            RIGHT_15_5: value  <= 0.34670698642730707340;
            RIGHT_15_6: value  <= 0.32944920659065252133;
            RIGHT_15_7: value  <= 0.38520970940589910336;
            RIGHT_15_8: value  <= 0.61500579118728637695;
            RIGHT_15_9: value  <= 0.53242927789688110352;
            RIGHT_15_10: value  <= 0.38430300354957580566;
            RIGHT_15_11: value  <= 0.57555872201919555664;
            RIGHT_15_12: value  <= 0.54714661836624145508;
            RIGHT_15_13: value  <= 0.61115288734436035156;
            RIGHT_15_14: value  <= 0.51895380020141601562;
            RIGHT_15_15: value  <= 0.47264769673347467593;
            RIGHT_15_16: value  <= 0.52603179216384887695;
            RIGHT_15_17: value  <= 0.39201408624649047852;
            RIGHT_15_18: value  <= 0.61196178197860717773;
            RIGHT_15_19: value  <= 0.53402662277221679688;
            RIGHT_15_20: value  <= 0.44551450014114379883;
            RIGHT_15_21: value  <= 0.53418618440628051758;
            RIGHT_15_22: value  <= 0.33616539835929870605;
            RIGHT_15_23: value  <= 0.08116444945335389571;
            RIGHT_15_24: value  <= 0.51898312568664550781;
            RIGHT_15_25: value  <= 0.23349590599536901303;
            RIGHT_15_26: value  <= 0.42956221103668207340;
            RIGHT_15_27: value  <= 0.55640292167663574219;
            RIGHT_15_28: value  <= 0.65791881084442138672;
            RIGHT_15_29: value  <= 0.36738881468772888184;
            RIGHT_15_30: value  <= 0.46421670913696289062;
            RIGHT_15_31: value  <= 0.27058771252632141113;
            RIGHT_15_32: value  <= 0.24490830302238458804;
            RIGHT_15_33: value  <= 0.55486911535263061523;
            RIGHT_15_34: value  <= 0.41036531329154968262;
            RIGHT_15_35: value  <= 0.48698890209197998047;
            RIGHT_15_36: value  <= 0.52876931428909301758;
            RIGHT_15_37: value  <= 0.46160620450973510742;
            RIGHT_15_38: value  <= 0.18198239803314208984;
            RIGHT_15_39: value  <= 0.52327787876129150391;
            RIGHT_15_40: value  <= 0.61765491962432861328;
            RIGHT_15_41: value  <= 0.43006989359855651855;
            RIGHT_15_42: value  <= 0.50008672475814819336;
            RIGHT_15_43: value  <= 0.67192137241363525391;
            RIGHT_15_44: value  <= 0.51781648397445678711;
            RIGHT_15_45: value  <= 0.62163108587265014648;
            RIGHT_15_46: value  <= 0.44100850820541381836;
            RIGHT_15_47: value  <= 0.54657220840454101562;
            RIGHT_15_48: value  <= 0.49958360195159912109;
            RIGHT_15_49: value  <= 0.52742338180541992188;
            RIGHT_15_50: value  <= 0.45722800493240361996;
            RIGHT_15_51: value  <= 0.41556000709533691406;
            RIGHT_15_52: value  <= 0.43530249595642089844;
            RIGHT_15_53: value  <= 0.67497581243515014648;
            RIGHT_15_54: value  <= 0.18832489848136899080;
            RIGHT_15_55: value  <= 0.52601581811904907227;
            RIGHT_15_56: value  <= 0.27764698863029479980;
            RIGHT_15_57: value  <= 0.46933171153068542480;
            RIGHT_15_58: value  <= 0.51697772741317749023;
            RIGHT_15_59: value  <= 0.51834410429000854492;
            RIGHT_15_60: value  <= 0.53621500730514526367;
            RIGHT_15_61: value  <= 0.43745940923690801450;
            RIGHT_15_62: value  <= 0.42093759775161737613;
            RIGHT_15_63: value  <= 0.47482660412788391113;
            RIGHT_15_64: value  <= 0.34245771169662481137;
            RIGHT_15_65: value  <= 0.63312637805938720703;
            RIGHT_15_66: value  <= 0.42268699407577520200;
            RIGHT_15_67: value  <= 0.54307800531387329102;
            RIGHT_15_68: value  <= 0.46976050734519958496;
            RIGHT_15_69: value  <= 0.53996050357818603516;
            RIGHT_15_70: value  <= 0.47473520040512090512;
            RIGHT_15_71: value  <= 0.55771100521087646484;
            RIGHT_15_72: value  <= 0.70239442586898803711;
            RIGHT_15_73: value  <= 0.38125100731849670410;
            RIGHT_15_74: value  <= 0.16878280043601989746;
            RIGHT_15_75: value  <= 0.63695681095123291016;
            RIGHT_15_76: value  <= 0.44876679778099060059;
            RIGHT_15_77: value  <= 0.29905700683593750000;
            RIGHT_15_78: value  <= 0.50784897804260253906;
            RIGHT_15_79: value  <= 0.52568262815475463867;
            RIGHT_15_80: value  <= 0.44942960143089288882;
            RIGHT_15_81: value  <= 0.26589488983154302426;
            RIGHT_15_82: value  <= 0.70872569084167480469;
            RIGHT_15_83: value  <= 0.37585180997848510742;
            RIGHT_15_84: value  <= 0.52385509014129638672;
            RIGHT_15_85: value  <= 0.58042472600936889648;
            RIGHT_15_86: value  <= 0.38730698823928827457;
            RIGHT_15_87: value  <= 0.56812518835067749023;
            RIGHT_15_88: value  <= 0.43182510137557977847;
            RIGHT_15_89: value  <= 0.43435549736022949219;
            RIGHT_15_90: value  <= 0.45375239849090581723;
            RIGHT_15_91: value  <= 0.41380101442337041684;
            RIGHT_15_92: value  <= 0.57171887159347534180;
            RIGHT_15_93: value  <= 0.52161228656768798828;
            RIGHT_15_94: value  <= 0.38183969259262090512;
            RIGHT_15_95: value  <= 0.42414000630378717593;
            RIGHT_15_96: value  <= 0.41869771480560302734;
            RIGHT_15_97: value  <= 0.52264511585235595703;
            RIGHT_15_98: value  <= 0.47157171368598937988;
            RIGHT_15_99: value  <= 0.33156448602676391602;
            RIGHT_15_100: value  <= 0.44581368565559392758;
            RIGHT_15_101: value  <= 0.36478888988494867496;
            RIGHT_15_102: value  <= 0.15679509937763211336;
            RIGHT_15_103: value  <= 0.62872701883316040039;
            RIGHT_15_104: value  <= 0.39437520503997802734;
            RIGHT_15_105: value  <= 0.50131380558013916016;
            RIGHT_15_106: value  <= 0.51287931203842163086;
            RIGHT_15_107: value  <= 0.57552158832550048828;
            RIGHT_15_108: value  <= 0.45580768585205078125;
            RIGHT_15_109: value  <= 0.21852590143680569734;
            RIGHT_15_110: value  <= 0.20906220376491549406;
            RIGHT_15_111: value  <= 0.71085482835769653320;
            RIGHT_15_112: value  <= 0.51561951637268066406;
            RIGHT_15_113: value  <= 0.44394320249557500668;
            RIGHT_15_114: value  <= 0.46204420924186712094;
            RIGHT_15_115: value  <= 0.54488998651504516602;
            RIGHT_15_116: value  <= 0.51336771249771118164;
            RIGHT_15_117: value  <= 0.64069348573684692383;
            RIGHT_15_118: value  <= 0.50155621767044067383;
            RIGHT_15_119: value  <= 0.51743787527084350586;
            RIGHT_15_120: value  <= 0.46778729557991027832;
            RIGHT_15_121: value  <= 0.10380929708480840512;
            RIGHT_15_122: value  <= 0.55320608615875244141;
            RIGHT_15_123: value  <= 0.52763891220092773438;
            RIGHT_15_124: value  <= 0.39320349693298339844;
            RIGHT_15_125: value  <= 0.47570338845252990723;
            RIGHT_15_126: value  <= 0.55357027053833007812;
            RIGHT_15_127: value  <= 0.51930642127990722656;
            RIGHT_15_128: value  <= 0.55936211347579956055;
            RIGHT_15_129: value  <= 0.47059568762779241391;
            RIGHT_15_130: value  <= 0.38100790977478027344;
            RIGHT_15_131: value  <= 0.61307388544082641602;
            RIGHT_15_132: value  <= 0.54293632507324218750;
            RIGHT_15_133: value  <= 0.41910758614540100098;
            RIGHT_15_134: value  <= 0.44716599583625787906;
            RIGHT_15_135: value  <= 0.46950098872184747867;
            RIGHT_15_136: value  <= 0.39458298683166498355;
            RIGHT_16_0: value  <= 0.38733118772506708316;
            RIGHT_16_1: value  <= 0.59739977121353149414;
            RIGHT_16_2: value  <= 0.25488111376762390137;
            RIGHT_16_3: value  <= 0.53872537612915039062;
            RIGHT_16_4: value  <= 0.35286578536033630371;
            RIGHT_16_5: value  <= 0.57659381628036499023;
            RIGHT_16_6: value  <= 0.55349981784820556641;
            RIGHT_16_7: value  <= 0.55478000640869140625;
            RIGHT_16_8: value  <= 0.45792970061302190610;
            RIGHT_16_9: value  <= 0.39040699601173400879;
            RIGHT_16_10: value  <= 0.52678012847900390625;
            RIGHT_16_11: value  <= 0.37143889069557189941;
            RIGHT_16_12: value  <= 0.41135668754577642270;
            RIGHT_16_13: value  <= 0.53293561935424804688;
            RIGHT_16_14: value  <= 0.37632051110267639160;
            RIGHT_16_15: value  <= 0.47052991390228271484;
            RIGHT_16_16: value  <= 0.55637162923812866211;
            RIGHT_16_17: value  <= 0.52151167392730712891;
            RIGHT_16_18: value  <= 0.30639201402664190121;
            RIGHT_16_19: value  <= 0.28859630227088928223;
            RIGHT_16_20: value  <= 0.58521968126296997070;
            RIGHT_16_21: value  <= 0.28700059652328491211;
            RIGHT_16_22: value  <= 0.46473708748817438297;
            RIGHT_16_23: value  <= 0.52470117807388305664;
            RIGHT_16_24: value  <= 0.59316617250442504883;
            RIGHT_16_25: value  <= 0.31303191184997558594;
            RIGHT_16_26: value  <= 0.50840771198272705078;
            RIGHT_16_27: value  <= 0.37407240271568298340;
            RIGHT_16_28: value  <= 0.74357217550277709961;
            RIGHT_16_29: value  <= 0.52805382013320922852;
            RIGHT_16_30: value  <= 0.34835430979728698730;
            RIGHT_16_31: value  <= 0.49323600530624389648;
            RIGHT_16_32: value  <= 0.22530519962310791016;
            RIGHT_16_33: value  <= 0.52646797895431518555;
            RIGHT_16_34: value  <= 0.70729321241378784180;
            RIGHT_16_35: value  <= 0.56682378053665161133;
            RIGHT_16_36: value  <= 0.57221567630767822266;
            RIGHT_16_37: value  <= 0.31146219372749328613;
            RIGHT_16_38: value  <= 0.52694618701934814453;
            RIGHT_16_39: value  <= 0.52457910776138305664;
            RIGHT_16_40: value  <= 0.46937671303749078922;
            RIGHT_16_41: value  <= 0.54090857505798339844;
            RIGHT_16_42: value  <= 0.44176620244979858398;
            RIGHT_16_43: value  <= 0.39734530448913568668;
            RIGHT_16_44: value  <= 0.52647268772125244141;
            RIGHT_16_45: value  <= 0.47498199343681341000;
            RIGHT_16_46: value  <= 0.33612239360809331723;
            RIGHT_16_47: value  <= 0.11726350337266920609;
            RIGHT_16_48: value  <= 0.13932949304580691252;
            RIGHT_16_49: value  <= 0.49211961030960077457;
            RIGHT_16_50: value  <= 0.50497019290924072266;
            RIGHT_16_51: value  <= 0.60487258434295654297;
            RIGHT_16_52: value  <= 0.46021929383277887515;
            RIGHT_16_53: value  <= 0.52260792255401611328;
            RIGHT_16_54: value  <= 0.33759570121765142270;
            RIGHT_16_55: value  <= 0.53035670518875122070;
            RIGHT_16_56: value  <= 0.39724540710449218750;
            RIGHT_16_57: value  <= 0.40634119510650640317;
            RIGHT_16_58: value  <= 0.68890458345413208008;
            RIGHT_16_59: value  <= 0.36247238516807561703;
            RIGHT_16_60: value  <= 0.50002872943878173828;
            RIGHT_16_61: value  <= 0.20028080046176910400;
            RIGHT_16_62: value  <= 0.63665360212326049805;
            RIGHT_16_63: value  <= 0.48678609728813171387;
            RIGHT_16_64: value  <= 0.53157979249954223633;
            RIGHT_16_65: value  <= 0.56052798032760620117;
            RIGHT_16_66: value  <= 0.51201480627059936523;
            RIGHT_16_67: value  <= 0.52073061466217041016;
            RIGHT_16_68: value  <= 0.46085759997367858887;
            RIGHT_16_69: value  <= 0.52422660589218139648;
            RIGHT_16_70: value  <= 0.37803208827972412109;
            RIGHT_16_71: value  <= 0.46118900179862981625;
            RIGHT_16_72: value  <= 0.58460158109664916992;
            RIGHT_16_73: value  <= 0.41845908761024480649;
            RIGHT_16_74: value  <= 0.52345657348632812500;
            RIGHT_16_75: value  <= 0.53564780950546264648;
            RIGHT_16_76: value  <= 0.23775640130043029785;
            RIGHT_16_77: value  <= 0.50504350662231445312;
            RIGHT_16_78: value  <= 0.46781000494956970215;
            RIGHT_16_79: value  <= 0.53236269950866699219;
            RIGHT_16_80: value  <= 0.56800121068954467773;
            RIGHT_16_81: value  <= 0.52968120574951171875;
            RIGHT_16_82: value  <= 0.74626070261001586914;
            RIGHT_16_83: value  <= 0.47521349787712102719;
            RIGHT_16_84: value  <= 0.50152552127838134766;
            RIGHT_16_85: value  <= 0.48962008953094482422;
            RIGHT_16_86: value  <= 0.53449410200119018555;
            RIGHT_16_87: value  <= 0.48039558529853820801;
            RIGHT_16_88: value  <= 0.76236087083816528320;
            RIGHT_16_89: value  <= 0.41916438937187200375;
            RIGHT_16_90: value  <= 0.53998219966888427734;
            RIGHT_16_91: value  <= 0.54249238967895507812;
            RIGHT_16_92: value  <= 0.45504111051559448242;
            RIGHT_16_93: value  <= 0.51891797780990600586;
            RIGHT_16_94: value  <= 0.47497498989105230160;
            RIGHT_16_95: value  <= 0.51775997877120971680;
            RIGHT_16_96: value  <= 0.51447242498397827148;
            RIGHT_16_97: value  <= 0.46673199534416198730;
            RIGHT_16_98: value  <= 0.61376398801803588867;
            RIGHT_16_99: value  <= 0.51935559511184692383;
            RIGHT_16_100: value  <= 0.30457559227943420410;
            RIGHT_16_101: value  <= 0.68875008821487426758;
            RIGHT_16_102: value  <= 0.50175631046295166016;
            RIGHT_16_103: value  <= 0.52426332235336303711;
            RIGHT_16_104: value  <= 0.47360289096832280942;
            RIGHT_16_105: value  <= 0.23898629844188690186;
            RIGHT_16_106: value  <= 0.44339430332183837891;
            RIGHT_16_107: value  <= 0.41488361358642578125;
            RIGHT_16_108: value  <= 0.06106159836053849654;
            RIGHT_16_109: value  <= 0.54238891601562500000;
            RIGHT_16_110: value  <= 0.53009921312332153320;
            RIGHT_16_111: value  <= 0.49573341012001037598;
            RIGHT_16_112: value  <= 0.28666600584983831235;
            RIGHT_16_113: value  <= 0.63181710243225097656;
            RIGHT_16_114: value  <= 0.49809598922729492188;
            RIGHT_16_115: value  <= 0.47080421447753911801;
            RIGHT_16_116: value  <= 0.49790981411933898926;
            RIGHT_16_117: value  <= 0.53779977560043334961;
            RIGHT_16_118: value  <= 0.55341911315917968750;
            RIGHT_16_119: value  <= 0.48252159357070917300;
            RIGHT_16_120: value  <= 0.40381389856338500977;
            RIGHT_16_121: value  <= 0.52600151300430297852;
            RIGHT_16_122: value  <= 0.76821839809417724609;
            RIGHT_16_123: value  <= 0.30622220039367681332;
            RIGHT_16_124: value  <= 0.46958100795745849609;
            RIGHT_16_125: value  <= 0.43869531154632568359;
            RIGHT_16_126: value  <= 0.58956301212310791016;
            RIGHT_16_127: value  <= 0.49424138665199279785;
            RIGHT_16_128: value  <= 0.45082521438598627261;
            RIGHT_16_129: value  <= 0.52238482236862182617;
            RIGHT_16_130: value  <= 0.35633018612861627750;
            RIGHT_16_131: value  <= 0.52188140153884887695;
            RIGHT_16_132: value  <= 0.51244372129440307617;
            RIGHT_16_133: value  <= 0.49197259545326227359;
            RIGHT_16_134: value  <= 0.46178871393203740903;
            RIGHT_16_135: value  <= 0.17127640545368200131;
            RIGHT_16_136: value  <= 0.51313877105712890625;
            RIGHT_16_137: value  <= 0.49979418516159057617;
            RIGHT_16_138: value  <= 0.55823111534118652344;
            RIGHT_16_139: value  <= 0.54524201154708862305;
            RIGHT_17_0: value  <= 0.59464621543884277344;
            RIGHT_17_1: value  <= 0.55778688192367553711;
            RIGHT_17_2: value  <= 0.32915300130844121762;
            RIGHT_17_3: value  <= 0.55459791421890258789;
            RIGHT_17_4: value  <= 0.55761402845382690430;
            RIGHT_17_5: value  <= 0.56453210115432739258;
            RIGHT_17_6: value  <= 0.70236331224441528320;
            RIGHT_17_7: value  <= 0.52892577648162841797;
            RIGHT_17_8: value  <= 0.40370491147041320801;
            RIGHT_17_9: value  <= 0.35578748583793640137;
            RIGHT_17_10: value  <= 0.46255499124526977539;
            RIGHT_17_11: value  <= 0.38696730136871337891;
            RIGHT_17_12: value  <= 0.53209269046783447266;
            RIGHT_17_13: value  <= 0.53633230924606323242;
            RIGHT_17_14: value  <= 0.32657089829444890805;
            RIGHT_17_15: value  <= 0.47741401195526117496;
            RIGHT_17_16: value  <= 0.54579311609268188477;
            RIGHT_17_17: value  <= 0.47931781411170959473;
            RIGHT_17_18: value  <= 0.35296788811683660336;
            RIGHT_17_19: value  <= 0.53529578447341918945;
            RIGHT_17_20: value  <= 0.38871330022811889648;
            RIGHT_17_21: value  <= 0.52736037969589233398;
            RIGHT_17_22: value  <= 0.68497377634048461914;
            RIGHT_17_23: value  <= 0.07022009044885639539;
            RIGHT_17_24: value  <= 0.51526021957397460938;
            RIGHT_17_25: value  <= 0.48972299695014948062;
            RIGHT_17_26: value  <= 0.38262099027633672543;
            RIGHT_17_27: value  <= 0.54219049215316772461;
            RIGHT_17_28: value  <= 0.50791162252426147461;
            RIGHT_17_29: value  <= 0.51284617185592651367;
            RIGHT_17_30: value  <= 0.43430820107460021973;
            RIGHT_17_31: value  <= 0.53599590063095092773;
            RIGHT_17_32: value  <= 0.51646977663040161133;
            RIGHT_17_33: value  <= 0.61140751838684082031;
            RIGHT_17_34: value  <= 0.50754940509796142578;
            RIGHT_17_35: value  <= 0.26887780427932739258;
            RIGHT_17_36: value  <= 0.67385399341583251953;
            RIGHT_17_37: value  <= 0.22127239406108858977;
            RIGHT_17_38: value  <= 0.45381900668144231625;
            RIGHT_17_39: value  <= 0.52474308013916015625;
            RIGHT_17_40: value  <= 0.39138820767402648926;
            RIGHT_17_41: value  <= 0.49902349710464477539;
            RIGHT_17_42: value  <= 0.50480902194976806641;
            RIGHT_17_43: value  <= 0.48423761129379272461;
            RIGHT_17_44: value  <= 0.25249770283699041196;
            RIGHT_17_45: value  <= 0.48984599113464361020;
            RIGHT_17_46: value  <= 0.22203169763088229094;
            RIGHT_17_47: value  <= 0.49338689446449279785;
            RIGHT_17_48: value  <= 0.37410449981689447574;
            RIGHT_17_49: value  <= 0.58180320262908935547;
            RIGHT_17_50: value  <= 0.52213358879089355469;
            RIGHT_17_51: value  <= 0.52312952280044555664;
            RIGHT_17_52: value  <= 0.47228169441223150082;
            RIGHT_17_53: value  <= 0.42424130439758300781;
            RIGHT_17_54: value  <= 0.56012850999832153320;
            RIGHT_17_55: value  <= 0.61366218328475952148;
            RIGHT_17_56: value  <= 0.45164099335670471191;
            RIGHT_17_57: value  <= 0.52949821949005126953;
            RIGHT_17_58: value  <= 0.52514511346817016602;
            RIGHT_17_59: value  <= 0.40655350685119628906;
            RIGHT_17_60: value  <= 0.49999570846557622739;
            RIGHT_17_61: value  <= 0.58134287595748901367;
            RIGHT_17_62: value  <= 0.55727928876876831055;
            RIGHT_17_63: value  <= 0.32128891348838811703;
            RIGHT_17_64: value  <= 0.45458820462226867676;
            RIGHT_17_65: value  <= 0.51522141695022583008;
            RIGHT_17_66: value  <= 0.37395030260086059570;
            RIGHT_17_67: value  <= 0.59382462501525878906;
            RIGHT_17_68: value  <= 0.41452041268348688297;
            RIGHT_17_69: value  <= 0.55149412155151367188;
            RIGHT_17_70: value  <= 0.46816679835319519043;
            RIGHT_17_71: value  <= 0.52291601896286010742;
            RIGHT_17_72: value  <= 0.36336138844490051270;
            RIGHT_17_73: value  <= 0.22117820382118230649;
            RIGHT_17_74: value  <= 0.57766091823577880859;
            RIGHT_17_75: value  <= 0.37566500902175897769;
            RIGHT_17_76: value  <= 0.56073749065399169922;
            RIGHT_17_77: value  <= 0.55182307958602905273;
            RIGHT_17_78: value  <= 0.59005767107009887695;
            RIGHT_17_79: value  <= 0.31563550233840942383;
            RIGHT_17_80: value  <= 0.58486622571945190430;
            RIGHT_17_81: value  <= 0.54836392402648925781;
            RIGHT_17_82: value  <= 0.37924841046333307437;
            RIGHT_17_83: value  <= 0.45769730210304260254;
            RIGHT_17_84: value  <= 0.56287872791290283203;
            RIGHT_17_85: value  <= 0.53910630941390991211;
            RIGHT_17_86: value  <= 0.47037428617477422543;
            RIGHT_17_87: value  <= 0.51918262243270874023;
            RIGHT_17_88: value  <= 0.34973978996276861020;
            RIGHT_17_89: value  <= 0.64083808660507202148;
            RIGHT_17_90: value  <= 0.52726852893829345703;
            RIGHT_17_91: value  <= 0.84165048599243164062;
            RIGHT_17_92: value  <= 0.43142348527908330746;
            RIGHT_17_93: value  <= 0.53825712203979492188;
            RIGHT_17_94: value  <= 0.47364759445190429688;
            RIGHT_17_95: value  <= 0.32815951108932500668;
            RIGHT_17_96: value  <= 0.51728862524032592773;
            RIGHT_17_97: value  <= 0.66876041889190673828;
            RIGHT_17_98: value  <= 0.47095969319343572446;
            RIGHT_17_99: value  <= 0.40598788857460021973;
            RIGHT_17_100: value  <= 0.66882789134979248047;
            RIGHT_17_101: value  <= 0.53442817926406860352;
            RIGHT_17_102: value  <= 0.16374860703945159912;
            RIGHT_17_103: value  <= 0.56332242488861083984;
            RIGHT_17_104: value  <= 0.47005268931388860532;
            RIGHT_17_105: value  <= 0.45361489057540888004;
            RIGHT_17_106: value  <= 0.44133889675140380859;
            RIGHT_17_107: value  <= 0.53564518690109252930;
            RIGHT_17_108: value  <= 0.37388110160827642270;
            RIGHT_17_109: value  <= 0.51888108253479003906;
            RIGHT_17_110: value  <= 0.55095332860946655273;
            RIGHT_17_111: value  <= 0.51954758167266845703;
            RIGHT_17_112: value  <= 0.45521140098571777344;
            RIGHT_17_113: value  <= 0.54974269866943359375;
            RIGHT_17_114: value  <= 0.54806441068649291992;
            RIGHT_17_115: value  <= 0.51785331964492797852;
            RIGHT_17_116: value  <= 0.57737642526626586914;
            RIGHT_17_117: value  <= 0.54608422517776489258;
            RIGHT_17_118: value  <= 0.52930849790573120117;
            RIGHT_17_119: value  <= 0.61219561100006103516;
            RIGHT_17_120: value  <= 0.51872807741165161133;
            RIGHT_17_121: value  <= 0.55761557817459106445;
            RIGHT_17_122: value  <= 0.50392812490463256836;
            RIGHT_17_123: value  <= 0.25258991122245788574;
            RIGHT_17_124: value  <= 0.54233711957931518555;
            RIGHT_17_125: value  <= 0.52130621671676635742;
            RIGHT_17_126: value  <= 0.42359098792076110840;
            RIGHT_17_127: value  <= 0.66240912675857543945;
            RIGHT_17_128: value  <= 0.40400519967079162598;
            RIGHT_17_129: value  <= 0.47951200604438781738;
            RIGHT_17_130: value  <= 0.53735041618347167969;
            RIGHT_17_131: value  <= 0.57593822479248046875;
            RIGHT_17_132: value  <= 0.35549798607826227359;
            RIGHT_17_133: value  <= 0.47317659854888921567;
            RIGHT_17_134: value  <= 0.70705670118331909180;
            RIGHT_17_135: value  <= 0.27817919850349431821;
            RIGHT_17_136: value  <= 0.50623041391372680664;
            RIGHT_17_137: value  <= 0.49345690011978149414;
            RIGHT_17_138: value  <= 0.34070080518722528629;
            RIGHT_17_139: value  <= 0.65790587663650512695;
            RIGHT_17_140: value  <= 0.50328421592712402344;
            RIGHT_17_141: value  <= 0.46950870752334600278;
            RIGHT_17_142: value  <= 0.51892018318176269531;
            RIGHT_17_143: value  <= 0.49401280283927917480;
            RIGHT_17_144: value  <= 0.45604279637336730957;
            RIGHT_17_145: value  <= 0.34839931130409240723;
            RIGHT_17_146: value  <= 0.50320827960968017578;
            RIGHT_17_147: value  <= 0.49149191379547119141;
            RIGHT_17_148: value  <= 0.56837642192840576172;
            RIGHT_17_149: value  <= 0.53334832191467285156;
            RIGHT_17_150: value  <= 0.43260601162910461426;
            RIGHT_17_151: value  <= 0.52015489339828491211;
            RIGHT_17_152: value  <= 0.49771949648857122250;
            RIGHT_17_153: value  <= 0.66669392585754394531;
            RIGHT_17_154: value  <= 0.42408201098442077637;
            RIGHT_17_155: value  <= 0.55638527870178222656;
            RIGHT_17_156: value  <= 0.47736850380897521973;
            RIGHT_17_157: value  <= 0.31712919473648071289;
            RIGHT_17_158: value  <= 0.70601707696914672852;
            RIGHT_17_159: value  <= 0.53307390213012695312;
            RIGHT_18_0: value  <= 0.68060368299484252930;
            RIGHT_18_1: value  <= 0.59657198190689086914;
            RIGHT_18_2: value  <= 0.34822869300842290707;
            RIGHT_18_3: value  <= 0.56933808326721191406;
            RIGHT_18_4: value  <= 0.54336887598037719727;
            RIGHT_18_5: value  <= 0.54843592643737792969;
            RIGHT_18_6: value  <= 0.54254651069641113281;
            RIGHT_18_7: value  <= 0.54295217990875244141;
            RIGHT_18_8: value  <= 0.53992640972137451172;
            RIGHT_18_9: value  <= 0.54402261972427368164;
            RIGHT_18_10: value  <= 0.54091197252273559570;
            RIGHT_18_11: value  <= 0.44790428876876831055;
            RIGHT_18_12: value  <= 0.57721698284149169922;
            RIGHT_18_13: value  <= 0.56858712434768676758;
            RIGHT_18_14: value  <= 0.52054089307785034180;
            RIGHT_18_15: value  <= 0.59806597232818603516;
            RIGHT_18_16: value  <= 0.29440331459045410156;
            RIGHT_18_17: value  <= 0.53771811723709106445;
            RIGHT_18_18: value  <= 0.52256888151168823242;
            RIGHT_18_19: value  <= 0.48923650383949279785;
            RIGHT_18_20: value  <= 0.56961381435394287109;
            RIGHT_18_21: value  <= 0.52256238460540771484;
            RIGHT_18_22: value  <= 0.46515759825706481934;
            RIGHT_18_23: value  <= 0.32863029837608337402;
            RIGHT_18_24: value  <= 0.50345462560653686523;
            RIGHT_18_25: value  <= 0.48890590667724609375;
            RIGHT_18_26: value  <= 0.38954809308052057437;
            RIGHT_18_27: value  <= 0.43724268674850458316;
            RIGHT_18_28: value  <= 0.50982052087783813477;
            RIGHT_18_29: value  <= 0.52465802431106567383;
            RIGHT_18_30: value  <= 0.39117100834846502133;
            RIGHT_18_31: value  <= 0.39427208900451660156;
            RIGHT_18_32: value  <= 0.50482118129730224609;
            RIGHT_18_33: value  <= 0.48726969957351690121;
            RIGHT_18_34: value  <= 0.62480747699737548828;
            RIGHT_18_35: value  <= 0.20000520348548889160;
            RIGHT_18_36: value  <= 0.53016197681427001953;
            RIGHT_18_37: value  <= 0.56531697511672973633;
            RIGHT_18_38: value  <= 0.50067067146301269531;
            RIGHT_18_39: value  <= 0.50463402271270751953;
            RIGHT_18_40: value  <= 0.47558510303497308902;
            RIGHT_18_41: value  <= 0.40046709775924682617;
            RIGHT_18_42: value  <= 0.49641749262809747867;
            RIGHT_18_43: value  <= 0.52180862426757812500;
            RIGHT_18_44: value  <= 0.53807932138442993164;
            RIGHT_18_45: value  <= 0.48774048686027532407;
            RIGHT_18_46: value  <= 0.36710259318351751157;
            RIGHT_18_47: value  <= 0.45790839195251470395;
            RIGHT_18_48: value  <= 0.51399451494216918945;
            RIGHT_18_49: value  <= 0.46642720699310302734;
            RIGHT_18_50: value  <= 0.51441830396652221680;
            RIGHT_18_51: value  <= 0.44140571355819702148;
            RIGHT_18_52: value  <= 0.61689937114715576172;
            RIGHT_18_53: value  <= 0.49748051166534418277;
            RIGHT_18_54: value  <= 0.39019080996513372250;
            RIGHT_18_55: value  <= 0.57904577255249023438;
            RIGHT_18_56: value  <= 0.50535911321640014648;
            RIGHT_18_57: value  <= 0.43298989534378051758;
            RIGHT_18_58: value  <= 0.66897618770599365234;
            RIGHT_18_59: value  <= 0.33778399229049682617;
            RIGHT_18_60: value  <= 0.53491330146789550781;
            RIGHT_18_61: value  <= 0.52282422780990600586;
            RIGHT_18_62: value  <= 0.42530721426010131836;
            RIGHT_18_63: value  <= 0.53789097070693969727;
            RIGHT_18_64: value  <= 0.47217491269111627750;
            RIGHT_18_65: value  <= 0.55483061075210571289;
            RIGHT_18_66: value  <= 0.42364639043807977847;
            RIGHT_18_67: value  <= 0.49693039059638982602;
            RIGHT_18_68: value  <= 0.16138119995594030209;
            RIGHT_18_69: value  <= 0.42230090498924260922;
            RIGHT_18_70: value  <= 0.60275578498840332031;
            RIGHT_18_71: value  <= 0.44224989414215087891;
            RIGHT_18_72: value  <= 0.66633248329162597656;
            RIGHT_18_73: value  <= 0.55269622802734375000;
            RIGHT_18_74: value  <= 0.33014988899230962582;
            RIGHT_18_75: value  <= 0.51750361919403076172;
            RIGHT_18_76: value  <= 0.53068768978118896484;
            RIGHT_18_77: value  <= 0.48365789651870727539;
            RIGHT_18_78: value  <= 0.51697367429733276367;
            RIGHT_18_79: value  <= 0.51639920473098754883;
            RIGHT_18_80: value  <= 0.37093898653984069824;
            RIGHT_18_81: value  <= 0.80539882183074951172;
            RIGHT_18_82: value  <= 0.46570208668708801270;
            RIGHT_18_83: value  <= 0.52587550878524780273;
            RIGHT_18_84: value  <= 0.38396438956260681152;
            RIGHT_18_85: value  <= 0.61870431900024414062;
            RIGHT_18_86: value  <= 0.49881500005722051450;
            RIGHT_18_87: value  <= 0.36320298910140991211;
            RIGHT_18_88: value  <= 0.57741481065750122070;
            RIGHT_18_89: value  <= 0.58582991361618041992;
            RIGHT_18_90: value  <= 0.50235372781753540039;
            RIGHT_18_91: value  <= 0.48537150025367742368;
            RIGHT_18_92: value  <= 0.36717799305915832520;
            RIGHT_18_93: value  <= 0.49946561455726617984;
            RIGHT_18_94: value  <= 0.62561017274856567383;
            RIGHT_18_95: value  <= 0.52818852663040161133;
            RIGHT_18_96: value  <= 0.55509579181671142578;
            RIGHT_18_97: value  <= 0.26133549213409418277;
            RIGHT_18_98: value  <= 0.50190317630767822266;
            RIGHT_18_99: value  <= 0.56616681814193725586;
            RIGHT_18_100: value  <= 0.55518132448196411133;
            RIGHT_18_101: value  <= 0.51513141393661499023;
            RIGHT_18_102: value  <= 0.44474598765373229980;
            RIGHT_18_103: value  <= 0.54878950119018554688;
            RIGHT_18_104: value  <= 0.51280808448791503906;
            RIGHT_18_105: value  <= 0.61015558242797851562;
            RIGHT_18_106: value  <= 0.41185480356216430664;
            RIGHT_18_107: value  <= 0.62523031234741210938;
            RIGHT_18_108: value  <= 0.36294108629226690121;
            RIGHT_18_109: value  <= 0.67380160093307495117;
            RIGHT_18_110: value  <= 0.52835988998413085938;
            RIGHT_18_111: value  <= 0.59007751941680908203;
            RIGHT_18_112: value  <= 0.60820537805557250977;
            RIGHT_18_113: value  <= 0.51809918880462646484;
            RIGHT_18_114: value  <= 0.40876251459121698550;
            RIGHT_18_115: value  <= 0.45385429263114929199;
            RIGHT_18_116: value  <= 0.41921341419219970703;
            RIGHT_18_117: value  <= 0.57062172889709472656;
            RIGHT_18_118: value  <= 0.58976382017135620117;
            RIGHT_18_119: value  <= 0.33576390147209167480;
            RIGHT_18_120: value  <= 0.13466019928455350008;
            RIGHT_18_121: value  <= 0.00061043637106195092;
            RIGHT_18_122: value  <= 0.70116281509399414062;
            RIGHT_18_123: value  <= 0.32828199863433837891;
            RIGHT_18_124: value  <= 0.45637390017509460449;
            RIGHT_18_125: value  <= 0.41039010882377630063;
            RIGHT_18_126: value  <= 0.54105907678604125977;
            RIGHT_18_127: value  <= 0.34382158517837518863;
            RIGHT_18_128: value  <= 0.44566130638122558594;
            RIGHT_18_129: value  <= 0.43626791238784790039;
            RIGHT_18_130: value  <= 0.65757977962493896484;
            RIGHT_18_131: value  <= 0.51373988389968872070;
            RIGHT_18_132: value  <= 0.49424308538436889648;
            RIGHT_18_133: value  <= 0.51175111532211303711;
            RIGHT_18_134: value  <= 0.25200259685516357422;
            RIGHT_18_135: value  <= 0.49278119206428527832;
            RIGHT_18_136: value  <= 0.36804521083831792660;
            RIGHT_18_137: value  <= 0.43636319041252141782;
            RIGHT_18_138: value  <= 0.45869469642639160156;
            RIGHT_18_139: value  <= 0.49204909801483148746;
            RIGHT_18_140: value  <= 0.49832528829574590512;
            RIGHT_18_141: value  <= 0.54900461435317993164;
            RIGHT_18_142: value  <= 0.50039529800415039062;
            RIGHT_18_143: value  <= 0.47215330600738530942;
            RIGHT_18_144: value  <= 0.49615910649299621582;
            RIGHT_18_145: value  <= 0.17410050332546231355;
            RIGHT_18_146: value  <= 0.47728818655014038086;
            RIGHT_18_147: value  <= 0.52927017211914062500;
            RIGHT_18_148: value  <= 0.40034240484237670898;
            RIGHT_18_149: value  <= 0.72129642963409423828;
            RIGHT_18_150: value  <= 0.55384761095046997070;
            RIGHT_18_151: value  <= 0.41632440686225891113;
            RIGHT_18_152: value  <= 0.45625001192092901059;
            RIGHT_18_153: value  <= 0.52802592515945434570;
            RIGHT_18_154: value  <= 0.52559971809387207031;
            RIGHT_18_155: value  <= 0.49520739912986760922;
            RIGHT_18_156: value  <= 0.55885308980941772461;
            RIGHT_18_157: value  <= 0.44238409399986272641;
            RIGHT_18_158: value  <= 0.52630358934402465820;
            RIGHT_18_159: value  <= 0.49984949827194208316;
            RIGHT_18_160: value  <= 0.48111200332641601562;
            RIGHT_18_161: value  <= 0.51769930124282836914;
            RIGHT_18_162: value  <= 0.54170542955398559570;
            RIGHT_18_163: value  <= 0.48940950632095342465;
            RIGHT_18_164: value  <= 0.45779189467430120297;
            RIGHT_18_165: value  <= 0.34004750847816467285;
            RIGHT_18_166: value  <= 0.50005030632019042969;
            RIGHT_18_167: value  <= 0.65975707769393920898;
            RIGHT_18_168: value  <= 0.49966529011726379395;
            RIGHT_18_169: value  <= 0.55037277936935424805;
            RIGHT_18_170: value  <= 0.52416700124740600586;
            RIGHT_18_171: value  <= 0.49744960665702819824;
            RIGHT_18_172: value  <= 0.58792287111282348633;
            RIGHT_18_173: value  <= 0.47052091360092157535;
            RIGHT_18_174: value  <= 0.37555369734764099121;
            RIGHT_18_175: value  <= 0.57907682657241821289;
            RIGHT_18_176: value  <= 0.39628401398658752441;
            RIGHT_19_0: value  <= 0.59619832038879394531;
            RIGHT_19_1: value  <= 0.44785520434379577637;
            RIGHT_19_2: value  <= 0.35782510042190551758;
            RIGHT_19_3: value  <= 0.30504280328750610352;
            RIGHT_19_4: value  <= 0.53446358442306518555;
            RIGHT_19_5: value  <= 0.55042648315429687500;
            RIGHT_19_6: value  <= 0.34760418534278869629;
            RIGHT_19_7: value  <= 0.62196469306945800781;
            RIGHT_19_8: value  <= 0.52780628204345703125;
            RIGHT_19_9: value  <= 0.37004441022872930356;
            RIGHT_19_10: value  <= 0.50919449329376220703;
            RIGHT_19_11: value  <= 0.54312258958816528320;
            RIGHT_19_12: value  <= 0.52213358879089355469;
            RIGHT_19_13: value  <= 0.47006508708000177554;
            RIGHT_19_14: value  <= 0.51409542560577392578;
            RIGHT_19_15: value  <= 0.48149210214614868164;
            RIGHT_19_16: value  <= 0.50258082151412963867;
            RIGHT_19_17: value  <= 0.68670457601547241211;
            RIGHT_19_18: value  <= 0.33506479859352111816;
            RIGHT_19_19: value  <= 0.52344137430191040039;
            RIGHT_19_20: value  <= 0.67225211858749389648;
            RIGHT_19_21: value  <= 0.27235329151153558902;
            RIGHT_19_22: value  <= 0.29069489240646362305;
            RIGHT_19_23: value  <= 0.63950210809707641602;
            RIGHT_19_24: value  <= 0.36566638946533197574;
            RIGHT_19_25: value  <= 0.47637018561363220215;
            RIGHT_19_26: value  <= 0.50309032201766967773;
            RIGHT_19_27: value  <= 0.51824611425399780273;
            RIGHT_19_28: value  <= 0.46949490904808038882;
            RIGHT_19_29: value  <= 0.42687839269638061523;
            RIGHT_19_30: value  <= 0.45716428756713872739;
            RIGHT_19_31: value  <= 0.32845470309257507324;
            RIGHT_19_32: value  <= 0.41793689131736760922;
            RIGHT_19_33: value  <= 0.53017157316207885742;
            RIGHT_19_34: value  <= 0.52207440137863159180;
            RIGHT_19_35: value  <= 0.41267579793930048160;
            RIGHT_19_36: value  <= 0.49945020675659179688;
            RIGHT_19_37: value  <= 0.49290320277214050293;
            RIGHT_19_38: value  <= 0.20398220419883730803;
            RIGHT_19_39: value  <= 0.57216948270797729492;
            RIGHT_19_40: value  <= 0.18018059432506561279;
            RIGHT_19_41: value  <= 0.48975929617881780453;
            RIGHT_19_42: value  <= 0.53837239742279052734;
            RIGHT_19_43: value  <= 0.57613271474838256836;
            RIGHT_19_44: value  <= 0.40976810455322271176;
            RIGHT_19_45: value  <= 0.50517761707305908203;
            RIGHT_19_46: value  <= 0.60318058729171752930;
            RIGHT_19_47: value  <= 0.54158830642700195312;
            RIGHT_19_48: value  <= 0.37022191286087041684;
            RIGHT_19_49: value  <= 0.48625651001930242368;
            RIGHT_19_50: value  <= 0.50889629125595092773;
            RIGHT_19_51: value  <= 0.61227089166641235352;
            RIGHT_19_52: value  <= 0.65561771392822265625;
            RIGHT_19_53: value  <= 0.16904720664024350252;
            RIGHT_19_54: value  <= 0.37252250313758850098;
            RIGHT_19_55: value  <= 0.49873429536819458008;
            RIGHT_19_56: value  <= 0.44648739695549011230;
            RIGHT_19_57: value  <= 0.34726628661155700684;
            RIGHT_19_58: value  <= 0.50048297643661499023;
            RIGHT_19_59: value  <= 0.45903238654136657715;
            RIGHT_19_60: value  <= 0.44970950484275817871;
            RIGHT_19_61: value  <= 0.42385208606719970703;
            RIGHT_19_62: value  <= 0.52581572532653808594;
            RIGHT_19_63: value  <= 0.54794532060623168945;
            RIGHT_19_64: value  <= 0.46746781468391418457;
            RIGHT_19_65: value  <= 0.55732029676437377930;
            RIGHT_19_66: value  <= 0.40741148591041570493;
            RIGHT_19_67: value  <= 0.58863520622253417969;
            RIGHT_19_68: value  <= 0.44871619343757629395;
            RIGHT_19_69: value  <= 0.28983271121978759766;
            RIGHT_19_70: value  <= 0.51978719234466552734;
            RIGHT_19_71: value  <= 0.49279558658599847965;
            RIGHT_19_72: value  <= 0.50125551223754882812;
            RIGHT_19_73: value  <= 0.56176078319549560547;
            RIGHT_19_74: value  <= 0.37655091285705571957;
            RIGHT_19_75: value  <= 0.48746308684349060059;
            RIGHT_19_76: value  <= 0.66913318634033203125;
            RIGHT_19_77: value  <= 0.27329459786415100098;
            RIGHT_19_78: value  <= 0.17820839583873748779;
            RIGHT_19_79: value  <= 0.32094758749008178711;
            RIGHT_19_80: value  <= 0.53072762489318847656;
            RIGHT_19_81: value  <= 0.51581299304962158203;
            RIGHT_19_82: value  <= 0.60755330324172973633;
            RIGHT_19_83: value  <= 0.52285957336425781250;
            RIGHT_19_84: value  <= 0.52156728506088256836;
            RIGHT_19_85: value  <= 0.43630391359329218082;
            RIGHT_19_86: value  <= 0.47898510098457341977;
            RIGHT_19_87: value  <= 0.53747731447219848633;
            RIGHT_19_88: value  <= 0.43661430478096008301;
            RIGHT_19_89: value  <= 0.58421492576599121094;
            RIGHT_19_90: value  <= 0.47210058569908142090;
            RIGHT_19_91: value  <= 0.43571090698242187500;
            RIGHT_19_92: value  <= 0.49918809533119201660;
            RIGHT_19_93: value  <= 0.49274989962577819824;
            RIGHT_19_94: value  <= 0.52458018064498901367;
            RIGHT_19_95: value  <= 0.57942241430282592773;
            RIGHT_19_96: value  <= 0.45445358753204351254;
            RIGHT_19_97: value  <= 0.55449050664901733398;
            RIGHT_19_98: value  <= 0.37802729010581970215;
            RIGHT_19_99: value  <= 0.48386740684509277344;
            RIGHT_19_100: value  <= 0.41636660695075988770;
            RIGHT_19_101: value  <= 0.53116250038146972656;
            RIGHT_19_102: value  <= 0.64665240049362182617;
            RIGHT_19_103: value  <= 0.21886579692363739014;
            RIGHT_19_104: value  <= 0.49588400125503540039;
            RIGHT_19_105: value  <= 0.46964588761329650879;
            RIGHT_19_106: value  <= 0.52171981334686279297;
            RIGHT_19_107: value  <= 0.48083150386810302734;
            RIGHT_19_108: value  <= 0.52282011508941650391;
            RIGHT_19_109: value  <= 0.57659977674484252930;
            RIGHT_19_110: value  <= 0.52531701326370239258;
            RIGHT_19_111: value  <= 0.17579819262027740479;
            RIGHT_19_112: value  <= 0.46949750185012817383;
            RIGHT_19_113: value  <= 0.33702209591865539551;
            RIGHT_19_114: value  <= 0.46945410966873168945;
            RIGHT_19_115: value  <= 0.27752599120140081235;
            RIGHT_19_116: value  <= 0.51926672458648681641;
            RIGHT_19_117: value  <= 0.61772608757019042969;
            RIGHT_19_118: value  <= 0.36847919225692749023;
            RIGHT_19_119: value  <= 0.48352020978927612305;
            RIGHT_19_120: value  <= 0.57230567932128906250;
            RIGHT_19_121: value  <= 0.52433192729949951172;
            RIGHT_19_122: value  <= 0.49687129259109502621;
            RIGHT_19_123: value  <= 0.43952131271362310239;
            RIGHT_19_124: value  <= 0.52698868513107299805;
            RIGHT_19_125: value  <= 0.50185042619705200195;
            RIGHT_19_126: value  <= 0.66983532905578613281;
            RIGHT_19_127: value  <= 0.53236472606658935547;
            RIGHT_19_128: value  <= 0.54398661851882934570;
            RIGHT_19_129: value  <= 0.55434262752532958984;
            RIGHT_19_130: value  <= 0.54267549514770507812;
            RIGHT_19_131: value  <= 0.35506111383438110352;
            RIGHT_19_132: value  <= 0.46306359767913818359;
            RIGHT_19_133: value  <= 0.55331951379776000977;
            RIGHT_19_134: value  <= 0.53224611282348632812;
            RIGHT_19_135: value  <= 0.54092890024185180664;
            RIGHT_19_136: value  <= 0.56288522481918334961;
            RIGHT_19_137: value  <= 0.27043169736862182617;
            RIGHT_19_138: value  <= 0.49805539846420288086;
            RIGHT_19_139: value  <= 0.50182962417602539062;
            RIGHT_19_140: value  <= 0.51852691173553466797;
            RIGHT_19_141: value  <= 0.56603360176086425781;
            RIGHT_19_142: value  <= 0.39571881294250488281;
            RIGHT_19_143: value  <= 0.50070542097091674805;
            RIGHT_19_144: value  <= 0.52284038066864013672;
            RIGHT_19_145: value  <= 0.59391832351684570312;
            RIGHT_19_146: value  <= 0.16333660483360290527;
            RIGHT_19_147: value  <= 0.49426248669624328613;
            RIGHT_19_148: value  <= 0.53287261724472045898;
            RIGHT_19_149: value  <= 0.49058890342712402344;
            RIGHT_19_150: value  <= 0.51380002498626708984;
            RIGHT_19_151: value  <= 0.50503468513488769531;
            RIGHT_19_152: value  <= 0.63778841495513916016;
            RIGHT_19_153: value  <= 0.41504821181297302246;
            RIGHT_19_154: value  <= 0.51497042179107666016;
            RIGHT_19_155: value  <= 0.48113578557968139648;
            RIGHT_19_156: value  <= 0.49923619627952581235;
            RIGHT_19_157: value  <= 0.48994860053062438965;
            RIGHT_19_158: value  <= 0.53926420211791992188;
            RIGHT_19_159: value  <= 0.37676128745079040527;
            RIGHT_19_160: value  <= 0.47479069232940668277;
            RIGHT_19_161: value  <= 0.54277169704437255859;
            RIGHT_19_162: value  <= 0.46186479926109308414;
            RIGHT_19_163: value  <= 0.48848950862884521484;
            RIGHT_19_164: value  <= 0.40171998739242548160;
            RIGHT_19_165: value  <= 0.26857739686965942383;
            RIGHT_19_166: value  <= 0.49797388911247247867;
            RIGHT_19_167: value  <= 0.55431222915649414062;
            RIGHT_19_168: value  <= 0.47099891304969787598;
            RIGHT_19_169: value  <= 0.53062361478805541992;
            RIGHT_19_170: value  <= 0.40517631173133850098;
            RIGHT_19_171: value  <= 0.47891938686370849609;
            RIGHT_19_172: value  <= 0.40118101239204412289;
            RIGHT_19_173: value  <= 0.50107032060623168945;
            RIGHT_19_174: value  <= 0.47731840610504150391;
            RIGHT_19_175: value  <= 0.51825290918350219727;
            RIGHT_19_176: value  <= 0.40981510281562810727;
            RIGHT_19_177: value  <= 0.54680430889129638672;
            RIGHT_19_178: value  <= 0.47838249802589422055;
            RIGHT_19_179: value  <= 0.52411228418350219727;
            RIGHT_19_180: value  <= 0.51136088371276855469;
            RIGHT_19_181: value  <= 0.54328018426895141602;
            RIGHT_20_0: value  <= 0.64211672544479370117;
            RIGHT_20_1: value  <= 0.67540389299392700195;
            RIGHT_20_2: value  <= 0.34233158826827997379;
            RIGHT_20_3: value  <= 0.54003179073333740234;
            RIGHT_20_4: value  <= 0.29350438714027410336;
            RIGHT_20_5: value  <= 0.53440642356872558594;
            RIGHT_20_6: value  <= 0.51320707798004150391;
            RIGHT_20_7: value  <= 0.55608451366424560547;
            RIGHT_20_8: value  <= 0.54047602415084838867;
            RIGHT_20_9: value  <= 0.55034661293029785156;
            RIGHT_20_10: value  <= 0.53697347640991210938;
            RIGHT_20_11: value  <= 0.52377498149871826172;
            RIGHT_20_12: value  <= 0.42235091328620910645;
            RIGHT_20_13: value  <= 0.47327259182929992676;
            RIGHT_20_14: value  <= 0.54327398538589477539;
            RIGHT_20_15: value  <= 0.60273271799087524414;
            RIGHT_20_16: value  <= 0.52139747142791748047;
            RIGHT_20_17: value  <= 0.47490629553794860840;
            RIGHT_20_18: value  <= 0.38434821367263788394;
            RIGHT_20_19: value  <= 0.34473359584808349609;
            RIGHT_20_20: value  <= 0.61939620971679687500;
            RIGHT_20_21: value  <= 0.53276282548904418945;
            RIGHT_20_22: value  <= 0.52749407291412353516;
            RIGHT_20_23: value  <= 0.49928390979766851254;
            RIGHT_20_24: value  <= 0.27666029334068298340;
            RIGHT_20_25: value  <= 0.52749711275100708008;
            RIGHT_20_26: value  <= 0.60011017322540283203;
            RIGHT_20_27: value  <= 0.52357178926467895508;
            RIGHT_20_28: value  <= 0.40343248844146728516;
            RIGHT_20_29: value  <= 0.45719841122627258301;
            RIGHT_20_30: value  <= 0.60346359014511108398;
            RIGHT_20_31: value  <= 0.53729712963104248047;
            RIGHT_20_32: value  <= 0.64378339052200317383;
            RIGHT_20_33: value  <= 0.53143328428268432617;
            RIGHT_20_34: value  <= 0.71308088302612304688;
            RIGHT_20_35: value  <= 0.53704041242599487305;
            RIGHT_20_36: value  <= 0.55144029855728149414;
            RIGHT_20_37: value  <= 0.59679841995239257812;
            RIGHT_20_38: value  <= 0.30185988545417791196;
            RIGHT_20_39: value  <= 0.44710969924926757812;
            RIGHT_20_40: value  <= 0.49899441003799438477;
            RIGHT_20_41: value  <= 0.50176489353179931641;
            RIGHT_20_42: value  <= 0.14820620417594909668;
            RIGHT_20_43: value  <= 0.59542238712310791016;
            RIGHT_20_44: value  <= 0.51960742473602294922;
            RIGHT_20_45: value  <= 0.48848581314086908511;
            RIGHT_20_46: value  <= 0.55788809061050415039;
            RIGHT_20_47: value  <= 0.53974777460098266602;
            RIGHT_20_48: value  <= 0.45332181453704828433;
            RIGHT_20_49: value  <= 0.42347279191017150879;
            RIGHT_20_50: value  <= 0.49584048986434942075;
            RIGHT_20_51: value  <= 0.71534800529479980469;
            RIGHT_20_52: value  <= 0.51949369907379150391;
            RIGHT_20_53: value  <= 0.60649001598358154297;
            RIGHT_20_54: value  <= 0.50608289241790771484;
            RIGHT_20_55: value  <= 0.52037787437438964844;
            RIGHT_20_56: value  <= 0.66269791126251220703;
            RIGHT_20_57: value  <= 0.35121849179267877750;
            RIGHT_20_58: value  <= 0.45298451185226440430;
            RIGHT_20_59: value  <= 0.53135812282562255859;
            RIGHT_20_60: value  <= 0.43333768844604492188;
            RIGHT_20_61: value  <= 0.40783908963203430176;
            RIGHT_20_62: value  <= 0.56438362598419189453;
            RIGHT_20_63: value  <= 0.52803301811218261719;
            RIGHT_20_64: value  <= 0.44077080488204961606;
            RIGHT_20_65: value  <= 0.24652279913425451108;
            RIGHT_20_66: value  <= 0.51396822929382324219;
            RIGHT_20_67: value  <= 0.59747868776321411133;
            RIGHT_20_68: value  <= 0.47687649726867681332;
            RIGHT_20_69: value  <= 0.52528268098831176758;
            RIGHT_20_70: value  <= 0.36295869946479797363;
            RIGHT_20_71: value  <= 0.43335610628128051758;
            RIGHT_20_72: value  <= 0.63310527801513671875;
            RIGHT_20_73: value  <= 0.45310580730438232422;
            RIGHT_20_74: value  <= 0.52571010589599609375;
            RIGHT_20_75: value  <= 0.45618548989295959473;
            RIGHT_20_76: value  <= 0.57369667291641235352;
            RIGHT_20_77: value  <= 0.45718750357627868652;
            RIGHT_20_78: value  <= 0.52201879024505615234;
            RIGHT_20_79: value  <= 0.52435082197189331055;
            RIGHT_20_80: value  <= 0.58990901708602905273;
            RIGHT_20_81: value  <= 0.28553789854049682617;
            RIGHT_20_82: value  <= 0.55064219236373901367;
            RIGHT_20_83: value  <= 0.51891750097274780273;
            RIGHT_20_84: value  <= 0.50407177209854125977;
            RIGHT_20_85: value  <= 0.48495069146156311035;
            RIGHT_20_86: value  <= 0.50320190191268920898;
            RIGHT_20_87: value  <= 0.58348792791366577148;
            RIGHT_20_88: value  <= 0.38964220881462102719;
            RIGHT_20_89: value  <= 0.52081221342086791992;
            RIGHT_20_90: value  <= 0.46412229537963872739;
            RIGHT_20_91: value  <= 0.43952199816703801938;
            RIGHT_20_92: value  <= 0.46810939908027648926;
            RIGHT_20_93: value  <= 0.40156200528144841977;
            RIGHT_20_94: value  <= 0.54528248310089111328;
            RIGHT_20_95: value  <= 0.48633798956871032715;
            RIGHT_20_96: value  <= 0.52474218606948852539;
            RIGHT_20_97: value  <= 0.36825248599052429199;
            RIGHT_20_98: value  <= 0.49612811207771301270;
            RIGHT_20_99: value  <= 0.48726621270179748535;
            RIGHT_20_100: value  <= 0.49509888887405401059;
            RIGHT_20_101: value  <= 0.53547459840774536133;
            RIGHT_20_102: value  <= 0.46388059854507451840;
            RIGHT_20_103: value  <= 0.46466401219367980957;
            RIGHT_20_104: value  <= 0.51302570104598999023;
            RIGHT_20_105: value  <= 0.56644618511199951172;
            RIGHT_20_106: value  <= 0.47158598899841308594;
            RIGHT_20_107: value  <= 0.30359649658203130551;
            RIGHT_20_108: value  <= 0.41070660948753362485;
            RIGHT_20_109: value  <= 0.49609071016311651059;
            RIGHT_20_110: value  <= 0.51409840583801269531;
            RIGHT_20_111: value  <= 0.62208187580108642578;
            RIGHT_20_112: value  <= 0.13224759697914120760;
            RIGHT_20_113: value  <= 0.50084167718887329102;
            RIGHT_20_114: value  <= 0.51301211118698120117;
            RIGHT_20_115: value  <= 0.49212029576301580258;
            RIGHT_20_116: value  <= 0.18591980636119839754;
            RIGHT_20_117: value  <= 0.55221217870712280273;
            RIGHT_20_118: value  <= 0.38564699888229370117;
            RIGHT_20_119: value  <= 0.54343092441558837891;
            RIGHT_20_120: value  <= 0.68406397104263305664;
            RIGHT_20_121: value  <= 0.53060990571975708008;
            RIGHT_20_122: value  <= 0.43781641125679021664;
            RIGHT_20_123: value  <= 0.06736146658658979935;
            RIGHT_20_124: value  <= 0.52556651830673217773;
            RIGHT_20_125: value  <= 0.44389671087265020200;
            RIGHT_20_126: value  <= 0.53995108604431152344;
            RIGHT_20_127: value  <= 0.50310248136520385742;
            RIGHT_20_128: value  <= 0.13983510434627530183;
            RIGHT_20_129: value  <= 0.49641060829162597656;
            RIGHT_20_130: value  <= 0.49463221430778497867;
            RIGHT_20_131: value  <= 0.52083408832550048828;
            RIGHT_20_132: value  <= 0.54261028766632080078;
            RIGHT_20_133: value  <= 0.51899671554565429688;
            RIGHT_20_134: value  <= 0.47521421313285827637;
            RIGHT_20_135: value  <= 0.63074797391891479492;
            RIGHT_20_136: value  <= 0.50268697738647460938;
            RIGHT_20_137: value  <= 0.38329708576202392578;
            RIGHT_20_138: value  <= 0.49698171019554138184;
            RIGHT_20_139: value  <= 0.69280272722244262695;
            RIGHT_20_140: value  <= 0.14764429628849029541;
            RIGHT_20_141: value  <= 0.48260560631752008609;
            RIGHT_20_142: value  <= 0.41296330094337457828;
            RIGHT_20_143: value  <= 0.37686121463775640317;
            RIGHT_20_144: value  <= 0.46374899148941040039;
            RIGHT_20_145: value  <= 0.53374791145324707031;
            RIGHT_20_146: value  <= 0.59003931283950805664;
            RIGHT_20_147: value  <= 0.43454289436340332031;
            RIGHT_20_148: value  <= 0.40513589978218078613;
            RIGHT_20_149: value  <= 0.55474412441253662109;
            RIGHT_20_150: value  <= 0.46725520491600042172;
            RIGHT_20_151: value  <= 0.50190007686614990234;
            RIGHT_20_152: value  <= 0.53636229038238525391;
            RIGHT_20_153: value  <= 0.57320207357406616211;
            RIGHT_20_154: value  <= 0.36350399255752557925;
            RIGHT_20_155: value  <= 0.45938020944595342465;
            RIGHT_20_156: value  <= 0.43391349911689758301;
            RIGHT_20_157: value  <= 0.54367768764495849609;
            RIGHT_20_158: value  <= 0.51762992143630981445;
            RIGHT_20_159: value  <= 0.56337797641754150391;
            RIGHT_20_160: value  <= 0.48008409142494201660;
            RIGHT_20_161: value  <= 0.51822227239608764648;
            RIGHT_20_162: value  <= 0.49357929825782781430;
            RIGHT_20_163: value  <= 0.53140252828598022461;
            RIGHT_20_164: value  <= 0.58962607383728027344;
            RIGHT_20_165: value  <= 0.50164777040481567383;
            RIGHT_20_166: value  <= 0.41268271207809448242;
            RIGHT_20_167: value  <= 0.58924478292465209961;
            RIGHT_20_168: value  <= 0.51894128322601318359;
            RIGHT_20_169: value  <= 0.49857059121131902524;
            RIGHT_20_170: value  <= 0.49558219313621520996;
            RIGHT_20_171: value  <= 0.50102657079696655273;
            RIGHT_20_172: value  <= 0.42263761162757867984;
            RIGHT_20_173: value  <= 0.58195871114730834961;
            RIGHT_20_174: value  <= 0.45117148756980901547;
            RIGHT_20_175: value  <= 0.51607340574264526367;
            RIGHT_20_176: value  <= 0.47361189126968378238;
            RIGHT_20_177: value  <= 0.33563950657844537906;
            RIGHT_20_178: value  <= 0.42640921473503107242;
            RIGHT_20_179: value  <= 0.57868278026580810547;
            RIGHT_20_180: value  <= 0.66778290271759033203;
            RIGHT_20_181: value  <= 0.43115469813346857242;
            RIGHT_20_182: value  <= 0.18888160586357119475;
            RIGHT_20_183: value  <= 0.58153688907623291016;
            RIGHT_20_184: value  <= 0.41325950622558588199;
            RIGHT_20_185: value  <= 0.48009279370307922363;
            RIGHT_20_186: value  <= 0.60414212942123413086;
            RIGHT_20_187: value  <= 0.30532771348953252621;
            RIGHT_20_188: value  <= 0.41788038611412048340;
            RIGHT_20_189: value  <= 0.48129200935363769531;
            RIGHT_20_190: value  <= 0.49717339873313898257;
            RIGHT_20_191: value  <= 0.52128481864929199219;
            RIGHT_20_192: value  <= 0.68920552730560302734;
            RIGHT_20_193: value  <= 0.43374860286712652035;
            RIGHT_20_194: value  <= 0.78437292575836181641;
            RIGHT_20_195: value  <= 0.53534239530563354492;
            RIGHT_20_196: value  <= 0.64259600639343261719;
            RIGHT_20_197: value  <= 0.51750177145004272461;
            RIGHT_20_198: value  <= 0.46289789676666259766;
            RIGHT_20_199: value  <= 0.32142710685729980469;
            RIGHT_20_200: value  <= 0.51416367292404174805;
            RIGHT_20_201: value  <= 0.63104897737503051758;
            RIGHT_20_202: value  <= 0.37232589721679687500;
            RIGHT_20_203: value  <= 0.48871129751205438785;
            RIGHT_20_204: value  <= 0.50039929151535034180;
            RIGHT_20_205: value  <= 0.56759268045425415039;
            RIGHT_20_206: value  <= 0.17772370576858520508;
            RIGHT_20_207: value  <= 0.54912507534027099609;
            RIGHT_20_208: value  <= 0.27907240390777587891;
            RIGHT_20_209: value  <= 0.49730318784713750668;
            RIGHT_20_210: value  <= 0.37767618894577031918;
            RIGHT_21_0: value  <= 0.40172868967056268863;
            RIGHT_21_1: value  <= 0.57464492321014404297;
            RIGHT_21_2: value  <= 0.55388098955154418945;
            RIGHT_21_3: value  <= 0.53826177120208740234;
            RIGHT_21_4: value  <= 0.55899268388748168945;
            RIGHT_21_5: value  <= 0.40203678607940668277;
            RIGHT_21_6: value  <= 0.33178439736366271973;
            RIGHT_21_7: value  <= 0.53079837560653686523;
            RIGHT_21_8: value  <= 0.64532989263534545898;
            RIGHT_21_9: value  <= 0.53705251216888427734;
            RIGHT_21_10: value  <= 0.38179719448089599609;
            RIGHT_21_11: value  <= 0.53820097446441650391;
            RIGHT_21_12: value  <= 0.55449652671813964844;
            RIGHT_21_13: value  <= 0.26788029074668878726;
            RIGHT_21_14: value  <= 0.52054339647293090820;
            RIGHT_21_15: value  <= 0.28613761067390441895;
            RIGHT_21_16: value  <= 0.52016979455947875977;
            RIGHT_21_17: value  <= 0.39598938822746282407;
            RIGHT_21_18: value  <= 0.52157157659530639648;
            RIGHT_21_19: value  <= 0.45844489336013788394;
            RIGHT_21_20: value  <= 0.53853511810302734375;
            RIGHT_21_21: value  <= 0.52935802936553955078;
            RIGHT_21_22: value  <= 0.50700891017913818359;
            RIGHT_21_23: value  <= 0.67264437675476074219;
            RIGHT_21_24: value  <= 0.55611097812652587891;
            RIGHT_21_25: value  <= 0.53086161613464355469;
            RIGHT_21_26: value  <= 0.46398720145225530453;
            RIGHT_21_27: value  <= 0.31418979167938232422;
            RIGHT_21_28: value  <= 0.53362947702407836914;
            RIGHT_21_29: value  <= 0.66034650802612304688;
            RIGHT_21_30: value  <= 0.45001828670501708984;
            RIGHT_21_31: value  <= 0.35997208952903747559;
            RIGHT_21_32: value  <= 0.49968141317367548160;
            RIGHT_21_33: value  <= 0.46847340464591979980;
            RIGHT_21_34: value  <= 0.18845909833908081055;
            RIGHT_21_35: value  <= 0.47990199923515319824;
            RIGHT_21_36: value  <= 0.35010111331939697266;
            RIGHT_21_37: value  <= 0.41176390647888178043;
            RIGHT_21_38: value  <= 0.53982460498809814453;
            RIGHT_21_39: value  <= 0.51791548728942871094;
            RIGHT_21_40: value  <= 0.23171770572662350740;
            RIGHT_21_41: value  <= 0.46436640620231628418;
            RIGHT_21_42: value  <= 0.44691911339759832211;
            RIGHT_21_43: value  <= 0.49259188771247858218;
            RIGHT_21_44: value  <= 0.39129018783569341489;
            RIGHT_21_45: value  <= 0.55017888545989990234;
            RIGHT_21_46: value  <= 0.46980848908424377441;
            RIGHT_21_47: value  <= 0.54808831214904785156;
            RIGHT_21_48: value  <= 0.50578862428665161133;
            RIGHT_21_49: value  <= 0.63982498645782470703;
            RIGHT_21_50: value  <= 0.62221372127532958984;
            RIGHT_21_51: value  <= 0.52221620082855224609;
            RIGHT_21_52: value  <= 0.49382260441780090332;
            RIGHT_21_53: value  <= 0.41167110204696660825;
            RIGHT_21_54: value  <= 0.46642690896987920590;
            RIGHT_21_55: value  <= 0.52497369050979614258;
            RIGHT_21_56: value  <= 0.50862592458724975586;
            RIGHT_21_57: value  <= 0.62034982442855834961;
            RIGHT_21_58: value  <= 0.50110971927642822266;
            RIGHT_21_59: value  <= 0.56283122301101684570;
            RIGHT_21_60: value  <= 0.46962749958038330078;
            RIGHT_21_61: value  <= 0.52876168489456176758;
            RIGHT_21_62: value  <= 0.50744771957397460938;
            RIGHT_21_63: value  <= 0.44896709918975830078;
            RIGHT_21_64: value  <= 0.52463638782501220703;
            RIGHT_21_65: value  <= 0.49051541090011602231;
            RIGHT_21_66: value  <= 0.64971512556076049805;
            RIGHT_21_67: value  <= 0.52276527881622314453;
            RIGHT_21_68: value  <= 0.38776180148124700375;
            RIGHT_21_69: value  <= 0.50238478183746337891;
            RIGHT_21_70: value  <= 0.54955857992172241211;
            RIGHT_21_71: value  <= 0.48595830798149108887;
            RIGHT_21_72: value  <= 0.43989309668540960141;
            RIGHT_21_73: value  <= 0.46050581336021417789;
            RIGHT_21_74: value  <= 0.29415771365165710449;
            RIGHT_21_75: value  <= 0.52185869216918945312;
            RIGHT_21_76: value  <= 0.54908162355422973633;
            RIGHT_21_77: value  <= 0.40813559293746948242;
            RIGHT_21_78: value  <= 0.52389502525329589844;
            RIGHT_21_79: value  <= 0.49080529808998107910;
            RIGHT_21_80: value  <= 0.52561181783676147461;
            RIGHT_21_81: value  <= 0.73136532306671142578;
            RIGHT_21_82: value  <= 0.45963698625564580746;
            RIGHT_21_83: value  <= 0.53088420629501342773;
            RIGHT_21_84: value  <= 0.45194861292839050293;
            RIGHT_21_85: value  <= 0.53607851266860961914;
            RIGHT_21_86: value  <= 0.54304420948028564453;
            RIGHT_21_87: value  <= 0.51460939645767211914;
            RIGHT_21_88: value  <= 0.18847459554672241211;
            RIGHT_21_89: value  <= 0.60938161611557006836;
            RIGHT_21_90: value  <= 0.46903759241104131528;
            RIGHT_21_91: value  <= 0.40460440516471857242;
            RIGHT_21_92: value  <= 0.52528482675552368164;
            RIGHT_21_93: value  <= 0.56901007890701293945;
            RIGHT_21_94: value  <= 0.17400950193405151367;
            RIGHT_21_95: value  <= 0.43548721075057977847;
            RIGHT_21_96: value  <= 0.43473169207572942563;
            RIGHT_21_97: value  <= 0.51605331897735595703;
            RIGHT_21_98: value  <= 0.72936528921127319336;
            RIGHT_21_99: value  <= 0.56331712007522583008;
            RIGHT_21_100: value  <= 0.51921367645263671875;
            RIGHT_21_101: value  <= 0.54179197549819946289;
            RIGHT_21_102: value  <= 0.52435618638992309570;
            RIGHT_21_103: value  <= 0.63870108127593994141;
            RIGHT_21_104: value  <= 0.29473468661308288574;
            RIGHT_21_105: value  <= 0.63088691234588623047;
            RIGHT_21_106: value  <= 0.42856499552726751157;
            RIGHT_21_107: value  <= 0.59415012598037719727;
            RIGHT_21_108: value  <= 0.58544808626174926758;
            RIGHT_21_109: value  <= 0.58490520715713500977;
            RIGHT_21_110: value  <= 0.52294230461120605469;
            RIGHT_21_111: value  <= 0.48983570933341979980;
            RIGHT_21_112: value  <= 0.54700392484664916992;
            RIGHT_21_113: value  <= 0.38429039716720581055;
            RIGHT_21_114: value  <= 0.28271919488906860352;
            RIGHT_21_115: value  <= 0.51488268375396728516;
            RIGHT_21_116: value  <= 0.70254462957382202148;
            RIGHT_21_117: value  <= 0.46560868620872497559;
            RIGHT_21_118: value  <= 0.51901197433471679688;
            RIGHT_21_119: value  <= 0.51617711782455444336;
            RIGHT_21_120: value  <= 0.46955159306526178531;
            RIGHT_21_121: value  <= 0.44258311390876770020;
            RIGHT_21_122: value  <= 0.42225030064582830258;
            RIGHT_21_123: value  <= 0.51799327135086059570;
            RIGHT_21_124: value  <= 0.76092642545700073242;
            RIGHT_21_125: value  <= 0.46717241406440740414;
            RIGHT_21_126: value  <= 0.14723660051822659578;
            RIGHT_21_127: value  <= 0.50165921449661254883;
            RIGHT_21_128: value  <= 0.56853622198104858398;
            RIGHT_21_129: value  <= 0.51379591226577758789;
            RIGHT_21_130: value  <= 0.37954080104827880859;
            RIGHT_21_131: value  <= 0.65804338455200195312;
            RIGHT_21_132: value  <= 0.40198868513107299805;
            RIGHT_21_133: value  <= 0.59544587135314941406;
            RIGHT_21_134: value  <= 0.51754468679428100586;
            RIGHT_21_135: value  <= 0.50571787357330322266;
            RIGHT_21_136: value  <= 0.80477148294448852539;
            RIGHT_21_137: value  <= 0.57199418544769287109;
            RIGHT_21_138: value  <= 0.49439039826393127441;
            RIGHT_21_139: value  <= 0.11433389782905580001;
            RIGHT_21_140: value  <= 0.56985741853713989258;
            RIGHT_21_141: value  <= 0.42187309265136718750;
            RIGHT_21_142: value  <= 0.46379259228706359863;
            RIGHT_21_143: value  <= 0.43820428848266601562;
            RIGHT_21_144: value  <= 0.51818847656250000000;
            RIGHT_21_145: value  <= 0.50893861055374145508;
            RIGHT_21_146: value  <= 0.50587952136993408203;
            RIGHT_21_147: value  <= 0.57930248975753784180;
            RIGHT_21_148: value  <= 0.53806531429290771484;
            RIGHT_21_149: value  <= 0.16847139596939089690;
            RIGHT_21_150: value  <= 0.67350268363952636719;
            RIGHT_21_151: value  <= 0.47757029533386230469;
            RIGHT_21_152: value  <= 0.23195350170135500822;
            RIGHT_21_153: value  <= 0.52629822492599487305;
            RIGHT_21_154: value  <= 0.35618188977241521664;
            RIGHT_21_155: value  <= 0.56190627813339233398;
            RIGHT_21_156: value  <= 0.67823082208633422852;
            RIGHT_21_157: value  <= 0.42907360196113591977;
            RIGHT_21_158: value  <= 0.55393511056900024414;
            RIGHT_21_159: value  <= 0.54341888427734375000;
            RIGHT_21_160: value  <= 0.65076571702957153320;
            RIGHT_21_161: value  <= 0.51617771387100219727;
            RIGHT_21_162: value  <= 0.42988368868827819824;
            RIGHT_21_163: value  <= 0.55824470520019531250;
            RIGHT_21_164: value  <= 0.07388007640838620271;
            RIGHT_21_165: value  <= 0.49775910377502441406;
            RIGHT_21_166: value  <= 0.54776942729949951172;
            RIGHT_21_167: value  <= 0.53133380413055419922;
            RIGHT_21_168: value  <= 0.53422421216964721680;
            RIGHT_21_169: value  <= 0.52044987678527832031;
            RIGHT_21_170: value  <= 0.41527429223060607910;
            RIGHT_21_171: value  <= 0.50188118219375610352;
            RIGHT_21_172: value  <= 0.35008639097213750668;
            RIGHT_21_173: value  <= 0.69686770439147949219;
            RIGHT_21_174: value  <= 0.50496298074722290039;
            RIGHT_21_175: value  <= 0.73211538791656494141;
            RIGHT_21_176: value  <= 0.51606708765029907227;
            RIGHT_21_177: value  <= 0.49497190117835998535;
            RIGHT_21_178: value  <= 0.45505958795547490903;
            RIGHT_21_179: value  <= 0.54435992240905761719;
            RIGHT_21_180: value  <= 0.38876569271087652035;
            RIGHT_21_181: value  <= 0.49717208743095397949;
            RIGHT_21_182: value  <= 0.50003677606582641602;
            RIGHT_21_183: value  <= 0.55603581666946411133;
            RIGHT_21_184: value  <= 0.46457770466804498843;
            RIGHT_21_185: value  <= 0.51934951543807983398;
            RIGHT_21_186: value  <= 0.34588789939880371094;
            RIGHT_21_187: value  <= 0.58701777458190917969;
            RIGHT_21_188: value  <= 0.53747731447219848633;
            RIGHT_21_189: value  <= 0.46409699320793151855;
            RIGHT_21_190: value  <= 0.67717897891998291016;
            RIGHT_21_191: value  <= 0.54280489683151245117;
            RIGHT_21_192: value  <= 0.46836739778518682309;
            RIGHT_21_193: value  <= 0.44242420792579650879;
            RIGHT_21_194: value  <= 0.51870870590209960938;
            RIGHT_21_195: value  <= 0.57712072134017944336;
            RIGHT_21_196: value  <= 0.56017017364501953125;
            RIGHT_21_197: value  <= 0.39147090911865228824;
            RIGHT_21_198: value  <= 0.56457388401031494141;
            RIGHT_21_199: value  <= 0.46927788853645330258;
            RIGHT_21_200: value  <= 0.37628141045570367984;
            RIGHT_21_201: value  <= 0.61515271663665771484;
            RIGHT_21_202: value  <= 0.43907511234283447266;
            RIGHT_21_203: value  <= 0.20630359649658200349;
            RIGHT_21_204: value  <= 0.51379072666168212891;
            RIGHT_21_205: value  <= 0.54275041818618774414;
            RIGHT_21_206: value  <= 0.47735071182250982114;
            RIGHT_21_207: value  <= 0.30349919199943542480;
            RIGHT_21_208: value  <= 0.44601860642433172055;
            RIGHT_21_209: value  <= 0.60274088382720947266;
            RIGHT_21_210: value  <= 0.51833057403564453125;
            RIGHT_21_211: value  <= 0.41887599229812622070;
            RIGHT_21_212: value  <= 0.65229612588882446289;

            default: value <= 0;

        endcase

    end

endmodule 
