module Feature_Threshold (

input int stage_num,
input int feature_num,
output real value

);

string name;
assign name = {"FEATURE_THRESH_", $sformatf("%d", stage_num), "_", $sformatf("%d", feature_num)};

always_comb
    begin

        case (name)

            "FEATURE_THRESH_0_0": value  <= 0.00401419587433338165;
            "FEATURE_THRESH_0_1": value  <= 0.01515133958309890054;
            "FEATURE_THRESH_0_2": value  <= 0.00421099318191409111;
            "FEATURE_THRESH_1_0": value  <= 0.00162271095905452967;
            "FEATURE_THRESH_1_1": value  <= 0.00229066493920981884;
            "FEATURE_THRESH_1_2": value  <= 0.00500257080420851707;
            "FEATURE_THRESH_1_3": value  <= 0.00796598941087722778;
            "FEATURE_THRESH_1_4": value  <= -0.00352270109578967094;
            "FEATURE_THRESH_1_5": value  <= 0.03666768968105320325;
            "FEATURE_THRESH_1_6": value  <= 0.00933614745736122131;
            "FEATURE_THRESH_1_7": value  <= 0.00869613140821456909;
            "FEATURE_THRESH_1_8": value  <= 0.00114888802636414766;
            "FEATURE_THRESH_1_9": value  <= -0.00214846897870302200;
            "FEATURE_THRESH_1_10": value  <= 0.00212190602906048298;
            "FEATURE_THRESH_1_11": value  <= -0.09394914656877520476;
            "FEATURE_THRESH_1_12": value  <= 0.00137777894269675016;
            "FEATURE_THRESH_1_13": value  <= 0.07306315749883650346;
            "FEATURE_THRESH_1_14": value  <= 0.00036767389974556863;
            "FEATURE_THRESH_1_15": value  <= -0.00604797108098864555;
            "FEATURE_THRESH_2_0": value  <= -0.01651068963110450052;
            "FEATURE_THRESH_2_1": value  <= 0.00270524993538856506;
            "FEATURE_THRESH_2_2": value  <= 0.00280698691494762897;
            "FEATURE_THRESH_2_3": value  <= -0.00154024001676589251;
            "FEATURE_THRESH_2_4": value  <= -0.00056386279175058007;
            "FEATURE_THRESH_2_5": value  <= 0.00192537298426032066;
            "FEATURE_THRESH_2_6": value  <= -0.00502148410305380821;
            "FEATURE_THRESH_2_7": value  <= 0.00263654207810759544;
            "FEATURE_THRESH_2_8": value  <= -0.00151277694385498762;
            "FEATURE_THRESH_2_9": value  <= -0.01015743985772129925;
            "FEATURE_THRESH_2_10": value  <= -0.01195366028696299987;
            "FEATURE_THRESH_2_11": value  <= 0.00488594919443130493;
            "FEATURE_THRESH_2_12": value  <= -0.08013291656970980559;
            "FEATURE_THRESH_2_13": value  <= 0.00106432801112532616;
            "FEATURE_THRESH_2_14": value  <= -0.00134194502606987953;
            "FEATURE_THRESH_2_15": value  <= -0.05460114032030109754;
            "FEATURE_THRESH_2_16": value  <= 0.00290716905146837234;
            "FEATURE_THRESH_2_17": value  <= 0.00074718717951327562;
            "FEATURE_THRESH_2_18": value  <= 0.00430138083174824715;
            "FEATURE_THRESH_2_19": value  <= 0.00450175721198320389;
            "FEATURE_THRESH_2_20": value  <= 0.02413850091397759870;
            "FEATURE_THRESH_3_0": value  <= 0.00192122301086783409;
            "FEATURE_THRESH_3_1": value  <= -0.00012748669541906565;
            "FEATURE_THRESH_3_2": value  <= 0.00051409931620582938;
            "FEATURE_THRESH_3_3": value  <= 0.00418786099180579185;
            "FEATURE_THRESH_3_4": value  <= 0.00510157179087400436;
            "FEATURE_THRESH_3_5": value  <= -0.00214484403841197491;
            "FEATURE_THRESH_3_6": value  <= -0.00289771193638443947;
            "FEATURE_THRESH_3_7": value  <= -0.02161067910492419850;
            "FEATURE_THRESH_3_8": value  <= -0.00462993187829852104;
            "FEATURE_THRESH_3_9": value  <= 0.00059393711853772402;
            "FEATURE_THRESH_3_10": value  <= 0.05387866124510769933;
            "FEATURE_THRESH_3_11": value  <= 0.00188873498700559139;
            "FEATURE_THRESH_3_12": value  <= -0.00236353394575417042;
            "FEATURE_THRESH_3_13": value  <= 0.02401779964566230080;
            "FEATURE_THRESH_3_14": value  <= 0.00020543030404951423;
            "FEATURE_THRESH_3_15": value  <= 0.00084790197433903813;
            "FEATURE_THRESH_3_16": value  <= 0.00140913296490907669;
            "FEATURE_THRESH_3_17": value  <= 0.00146426295395940542;
            "FEATURE_THRESH_3_18": value  <= 0.00163525494281202555;
            "FEATURE_THRESH_3_19": value  <= 0.00083172752056270838;
            "FEATURE_THRESH_3_20": value  <= -0.00209988909773528576;
            "FEATURE_THRESH_3_21": value  <= -0.00074213981861248612;
            "FEATURE_THRESH_3_22": value  <= 0.00326550495810806751;
            "FEATURE_THRESH_3_23": value  <= 0.00089134991867467761;
            "FEATURE_THRESH_3_24": value  <= -0.01528417970985170016;
            "FEATURE_THRESH_3_25": value  <= 0.00483814114704728127;
            "FEATURE_THRESH_3_26": value  <= -0.00091093179071322083;
            "FEATURE_THRESH_3_27": value  <= -0.00612750602886080742;
            "FEATURE_THRESH_3_28": value  <= -0.00044576259097084403;
            "FEATURE_THRESH_3_29": value  <= 0.02264654077589510137;
            "FEATURE_THRESH_3_30": value  <= -0.00188049604184925556;
            "FEATURE_THRESH_3_31": value  <= 0.00708891078829765320;
            "FEATURE_THRESH_3_32": value  <= 0.00173180503770709038;
            "FEATURE_THRESH_3_33": value  <= -0.00684827007353305817;
            "FEATURE_THRESH_3_34": value  <= -0.00001506253011029912;
            "FEATURE_THRESH_3_35": value  <= 0.02947556972503660028;
            "FEATURE_THRESH_3_36": value  <= 0.00813873298466205597;
            "FEATURE_THRESH_3_37": value  <= 0.02094295062124729850;
            "FEATURE_THRESH_3_38": value  <= -0.00956655293703079224;
            "FEATURE_THRESH_4_0": value  <= -0.00028206960996612906;
            "FEATURE_THRESH_4_1": value  <= 0.00167906004935503006;
            "FEATURE_THRESH_4_2": value  <= 0.00069827912375330925;
            "FEATURE_THRESH_4_3": value  <= 0.00078959012171253562;
            "FEATURE_THRESH_4_4": value  <= -0.00285604991950094700;
            "FEATURE_THRESH_4_5": value  <= -0.00381224695593118668;
            "FEATURE_THRESH_4_6": value  <= 0.00158966204617172480;
            "FEATURE_THRESH_4_7": value  <= 0.01007833983749150016;
            "FEATURE_THRESH_4_8": value  <= -0.06352630257606510511;
            "FEATURE_THRESH_4_9": value  <= -0.00910314917564392090;
            "FEATURE_THRESH_4_10": value  <= -0.00240350002422928810;
            "FEATURE_THRESH_4_11": value  <= 0.00152263604104518890;
            "FEATURE_THRESH_4_12": value  <= 0.01799743995070459887;
            "FEATURE_THRESH_4_13": value  <= -0.00645381910726428032;
            "FEATURE_THRESH_4_14": value  <= -0.01188076008111240041;
            "FEATURE_THRESH_4_15": value  <= 0.00127136602532118559;
            "FEATURE_THRESH_4_16": value  <= 0.00113761099055409431;
            "FEATURE_THRESH_4_17": value  <= -0.00426519988104701042;
            "FEATURE_THRESH_4_18": value  <= -0.00296028610318899155;
            "FEATURE_THRESH_4_19": value  <= -0.00884482264518737793;
            "FEATURE_THRESH_4_20": value  <= -0.00664306897670030594;
            "FEATURE_THRESH_4_21": value  <= 0.00399978086352348328;
            "FEATURE_THRESH_4_22": value  <= -0.00412217201665043831;
            "FEATURE_THRESH_4_23": value  <= 0.01562490966171030046;
            "FEATURE_THRESH_4_24": value  <= -0.01035641971975569987;
            "FEATURE_THRESH_4_25": value  <= -0.00879608094692230225;
            "FEATURE_THRESH_4_26": value  <= 0.16226939857006070222;
            "FEATURE_THRESH_4_27": value  <= 0.00455425307154655457;
            "FEATURE_THRESH_4_28": value  <= -0.00213092099875211716;
            "FEATURE_THRESH_4_29": value  <= -0.01320842001587150052;
            "FEATURE_THRESH_4_30": value  <= -0.06599667668342590332;
            "FEATURE_THRESH_4_31": value  <= 0.00791426561772823334;
            "FEATURE_THRESH_4_32": value  <= 0.02089427970349790054;
            "FEATURE_THRESH_5_0": value  <= 0.00119611597619950771;
            "FEATURE_THRESH_5_1": value  <= -0.00186798302456736565;
            "FEATURE_THRESH_5_2": value  <= -0.00019579799845814705;
            "FEATURE_THRESH_5_3": value  <= -0.00080255657667294145;
            "FEATURE_THRESH_5_4": value  <= -0.00245108106173574924;
            "FEATURE_THRESH_5_5": value  <= 0.00050361850298941135;
            "FEATURE_THRESH_5_6": value  <= 0.00402933498844504356;
            "FEATURE_THRESH_5_7": value  <= -0.01445170957595109940;
            "FEATURE_THRESH_5_8": value  <= 0.00203809794038534164;
            "FEATURE_THRESH_5_9": value  <= -0.00161551905330270529;
            "FEATURE_THRESH_5_10": value  <= 0.00334583409130573273;
            "FEATURE_THRESH_5_11": value  <= 0.00163795799016952515;
            "FEATURE_THRESH_5_12": value  <= 0.03025121055543419923;
            "FEATURE_THRESH_5_13": value  <= 0.03725199028849599664;
            "FEATURE_THRESH_5_14": value  <= -0.02510979026556019872;
            "FEATURE_THRESH_5_15": value  <= -0.00530990585684776306;
            "FEATURE_THRESH_5_16": value  <= 0.00120864796917885542;
            "FEATURE_THRESH_5_17": value  <= -0.02190767973661419954;
            "FEATURE_THRESH_5_18": value  <= 0.00541165797039866447;
            "FEATURE_THRESH_5_19": value  <= 0.06994632631540299850;
            "FEATURE_THRESH_5_20": value  <= 0.00034520021290518343;
            "FEATURE_THRESH_5_21": value  <= 0.00126277096569538116;
            "FEATURE_THRESH_5_22": value  <= 0.02271950989961619982;
            "FEATURE_THRESH_5_23": value  <= -0.00181110005360096693;
            "FEATURE_THRESH_5_24": value  <= 0.00334696704521775246;
            "FEATURE_THRESH_5_25": value  <= 0.00040791751234792173;
            "FEATURE_THRESH_5_26": value  <= 0.01273479964584110086;
            "FEATURE_THRESH_5_27": value  <= -0.00731197278946638107;
            "FEATURE_THRESH_5_28": value  <= -0.05694875121116640265;
            "FEATURE_THRESH_5_29": value  <= -0.00501165911555290222;
            "FEATURE_THRESH_5_30": value  <= 0.00603343686088919640;
            "FEATURE_THRESH_5_31": value  <= 0.00394374411553144455;
            "FEATURE_THRESH_5_32": value  <= -0.00365911191329360008;
            "FEATURE_THRESH_5_33": value  <= -0.00384561810642480850;
            "FEATURE_THRESH_5_34": value  <= -0.00719262612983584404;
            "FEATURE_THRESH_5_35": value  <= -0.05279894173145290026;
            "FEATURE_THRESH_5_36": value  <= -0.00795376673340797424;
            "FEATURE_THRESH_5_37": value  <= -0.00273441802710294724;
            "FEATURE_THRESH_5_38": value  <= -0.00185079395305365324;
            "FEATURE_THRESH_5_39": value  <= 0.01591891981661320080;
            "FEATURE_THRESH_5_40": value  <= -0.00126876798458397388;
            "FEATURE_THRESH_5_41": value  <= 0.00628839107230305672;
            "FEATURE_THRESH_5_42": value  <= -0.00622598920017480850;
            "FEATURE_THRESH_5_43": value  <= -0.01213259994983669973;
            "FEATURE_THRESH_6_0": value  <= -0.00391849083825945854;
            "FEATURE_THRESH_6_1": value  <= 0.00159712997265160084;
            "FEATURE_THRESH_6_2": value  <= 0.01778011023998260151;
            "FEATURE_THRESH_6_3": value  <= 0.00065334769897162914;
            "FEATURE_THRESH_6_4": value  <= -0.00028353091329336166;
            "FEATURE_THRESH_6_5": value  <= 0.00161046895664185286;
            "FEATURE_THRESH_6_6": value  <= -0.09775061905384059557;
            "FEATURE_THRESH_6_7": value  <= 0.00055182358482852578;
            "FEATURE_THRESH_6_8": value  <= -0.01285822037607430024;
            "FEATURE_THRESH_6_9": value  <= 0.00415302393957972527;
            "FEATURE_THRESH_6_10": value  <= 0.00170924596022814512;
            "FEATURE_THRESH_6_11": value  <= 0.00752173596993088722;
            "FEATURE_THRESH_6_12": value  <= 0.00224798102863132954;
            "FEATURE_THRESH_6_13": value  <= 0.05200621113181110033;
            "FEATURE_THRESH_6_14": value  <= 0.01208552997559310047;
            "FEATURE_THRESH_6_15": value  <= 0.00001468782011215808;
            "FEATURE_THRESH_6_16": value  <= 0.00000713951885700226;
            "FEATURE_THRESH_6_17": value  <= -0.00460016401484608650;
            "FEATURE_THRESH_6_18": value  <= 0.00200589490123093128;
            "FEATURE_THRESH_6_19": value  <= 0.00450502708554267883;
            "FEATURE_THRESH_6_20": value  <= 0.01174683030694720007;
            "FEATURE_THRESH_6_21": value  <= -0.05831633880734440195;
            "FEATURE_THRESH_6_22": value  <= 0.00023629379575140774;
            "FEATURE_THRESH_6_23": value  <= -0.00781561806797981262;
            "FEATURE_THRESH_6_24": value  <= -0.01087616011500359969;
            "FEATURE_THRESH_6_25": value  <= -0.00277455197647213936;
            "FEATURE_THRESH_6_26": value  <= -0.00078276381827890873;
            "FEATURE_THRESH_6_27": value  <= 0.01387040968984369974;
            "FEATURE_THRESH_6_28": value  <= -0.02367491088807580080;
            "FEATURE_THRESH_6_29": value  <= -0.00001487940971856006;
            "FEATURE_THRESH_6_30": value  <= 0.00361906411126255989;
            "FEATURE_THRESH_6_31": value  <= -0.01981711015105249926;
            "FEATURE_THRESH_6_32": value  <= -0.00381540390662848949;
            "FEATURE_THRESH_6_33": value  <= -0.00497758295387029648;
            "FEATURE_THRESH_6_34": value  <= 0.00224410207010805607;
            "FEATURE_THRESH_6_35": value  <= 0.01228245999664069957;
            "FEATURE_THRESH_6_36": value  <= -0.00285486993379890919;
            "FEATURE_THRESH_6_37": value  <= -0.00378756690770387650;
            "FEATURE_THRESH_6_38": value  <= -0.00122012302745133638;
            "FEATURE_THRESH_6_39": value  <= 0.01016059983521700079;
            "FEATURE_THRESH_6_40": value  <= -0.01617456972599029888;
            "FEATURE_THRESH_6_41": value  <= 0.01929246075451369891;
            "FEATURE_THRESH_6_42": value  <= -0.00324795395135879517;
            "FEATURE_THRESH_6_43": value  <= -0.00938034802675247192;
            "FEATURE_THRESH_6_44": value  <= -0.01260612998157739986;
            "FEATURE_THRESH_6_45": value  <= -0.02562193013727660090;
            "FEATURE_THRESH_6_46": value  <= -0.00007574149640277028;
            "FEATURE_THRESH_6_47": value  <= -0.08921088278293609619;
            "FEATURE_THRESH_6_48": value  <= -0.00276704807765781879;
            "FEATURE_THRESH_6_49": value  <= 0.00027152578695677221;
            "FEATURE_THRESH_7_0": value  <= 0.00147862196899950504;
            "FEATURE_THRESH_7_1": value  <= -0.00187416595872491598;
            "FEATURE_THRESH_7_2": value  <= -0.00171510095242410898;
            "FEATURE_THRESH_7_3": value  <= -0.00189392699394375086;
            "FEATURE_THRESH_7_4": value  <= -0.00530060520395636559;
            "FEATURE_THRESH_7_5": value  <= -0.04666253179311750238;
            "FEATURE_THRESH_7_6": value  <= -0.00079431332414969802;
            "FEATURE_THRESH_7_7": value  <= 0.01489167008548980022;
            "FEATURE_THRESH_7_8": value  <= -0.00120465294457972050;
            "FEATURE_THRESH_7_9": value  <= 0.00606193812564015388;
            "FEATURE_THRESH_7_10": value  <= -0.00252866488881409168;
            "FEATURE_THRESH_7_11": value  <= -0.00590102188289165497;
            "FEATURE_THRESH_7_12": value  <= 0.00567027600482106209;
            "FEATURE_THRESH_7_13": value  <= -0.00303041003644466400;
            "FEATURE_THRESH_7_14": value  <= 0.00298036495223641396;
            "FEATURE_THRESH_7_15": value  <= -0.07584051042795179887;
            "FEATURE_THRESH_7_16": value  <= 0.01926253922283650138;
            "FEATURE_THRESH_7_17": value  <= 0.00018888259364757687;
            "FEATURE_THRESH_7_18": value  <= 0.02936954982578749915;
            "FEATURE_THRESH_7_19": value  <= 0.00104176194872707129;
            "FEATURE_THRESH_7_20": value  <= 0.00261256401427090168;
            "FEATURE_THRESH_7_21": value  <= 0.00096977467183023691;
            "FEATURE_THRESH_7_22": value  <= 0.00059512659208849072;
            "FEATURE_THRESH_7_23": value  <= -0.10156559944152830643;
            "FEATURE_THRESH_7_24": value  <= 0.03615669906139370310;
            "FEATURE_THRESH_7_25": value  <= 0.00346241402439773083;
            "FEATURE_THRESH_7_26": value  <= 0.01955498009920119892;
            "FEATURE_THRESH_7_27": value  <= -0.00231214403174817562;
            "FEATURE_THRESH_7_28": value  <= -0.00186052895151078701;
            "FEATURE_THRESH_7_29": value  <= -0.00094026362057775259;
            "FEATURE_THRESH_7_30": value  <= -0.00524183316156268120;
            "FEATURE_THRESH_7_31": value  <= 0.00011729019752237946;
            "FEATURE_THRESH_7_32": value  <= 0.00118788401596248150;
            "FEATURE_THRESH_7_33": value  <= -0.01088135968893770046;
            "FEATURE_THRESH_7_34": value  <= 0.00173548597376793623;
            "FEATURE_THRESH_7_35": value  <= -0.00651190523058176041;
            "FEATURE_THRESH_7_36": value  <= -0.00121364300139248371;
            "FEATURE_THRESH_7_37": value  <= -0.01035424042493100077;
            "FEATURE_THRESH_7_38": value  <= 0.00055858830455690622;
            "FEATURE_THRESH_7_39": value  <= 0.01529964990913870032;
            "FEATURE_THRESH_7_40": value  <= -0.02158821001648900118;
            "FEATURE_THRESH_7_41": value  <= -0.12834629416465759277;
            "FEATURE_THRESH_7_42": value  <= -0.00229271897114813328;
            "FEATURE_THRESH_7_43": value  <= 0.07991510629653930664;
            "FEATURE_THRESH_7_44": value  <= -0.07944109290838240189;
            "FEATURE_THRESH_7_45": value  <= -0.00528000108897686005;
            "FEATURE_THRESH_7_46": value  <= 0.00104631099384278059;
            "FEATURE_THRESH_7_47": value  <= 0.00026317298761568964;
            "FEATURE_THRESH_7_48": value  <= -0.00361731601879000664;
            "FEATURE_THRESH_7_49": value  <= 0.01142187975347040002;
            "FEATURE_THRESH_7_50": value  <= -0.00199632789008319378;
            "FEATURE_THRESH_8_0": value  <= -0.00996912457048892975;
            "FEATURE_THRESH_8_1": value  <= 0.00073073059320449829;
            "FEATURE_THRESH_8_2": value  <= 0.00064045301405712962;
            "FEATURE_THRESH_8_3": value  <= 0.00454240199178457260;
            "FEATURE_THRESH_8_4": value  <= 0.00009247744310414420;
            "FEATURE_THRESH_8_5": value  <= -0.00866031460464000702;
            "FEATURE_THRESH_8_6": value  <= 0.00805158168077468872;
            "FEATURE_THRESH_8_7": value  <= 0.00043835240649059415;
            "FEATURE_THRESH_8_8": value  <= -0.00009816897363634781;
            "FEATURE_THRESH_8_9": value  <= -0.00112987903412431479;
            "FEATURE_THRESH_8_10": value  <= 0.00643561501055955887;
            "FEATURE_THRESH_8_11": value  <= -0.05682932958006860213;
            "FEATURE_THRESH_8_12": value  <= 0.00406681699678301811;
            "FEATURE_THRESH_8_13": value  <= 0.00004816479849978351;
            "FEATURE_THRESH_8_14": value  <= 0.00617950176820158958;
            "FEATURE_THRESH_8_15": value  <= 0.00649857521057128906;
            "FEATURE_THRESH_8_16": value  <= -0.00102110905572772026;
            "FEATURE_THRESH_8_17": value  <= -0.00542475283145904541;
            "FEATURE_THRESH_8_18": value  <= -0.00105598999653011560;
            "FEATURE_THRESH_8_19": value  <= 0.00066465808777138591;
            "FEATURE_THRESH_8_20": value  <= -0.00027524109464138746;
            "FEATURE_THRESH_8_21": value  <= 0.00422932021319866180;
            "FEATURE_THRESH_8_22": value  <= -0.00328682106919586658;
            "FEATURE_THRESH_8_23": value  <= 0.00015611879643984139;
            "FEATURE_THRESH_8_24": value  <= -0.00000736213814889197;
            "FEATURE_THRESH_8_25": value  <= -0.01476725004613400026;
            "FEATURE_THRESH_8_26": value  <= 0.02448959089815620077;
            "FEATURE_THRESH_8_27": value  <= -0.00037652091123163700;
            "FEATURE_THRESH_8_28": value  <= 0.00000736576885174145;
            "FEATURE_THRESH_8_29": value  <= -0.01509993989020590004;
            "FEATURE_THRESH_8_30": value  <= -0.00383166503161191940;
            "FEATURE_THRESH_8_31": value  <= 0.01692540012300009986;
            "FEATURE_THRESH_8_32": value  <= -0.00304778502322733402;
            "FEATURE_THRESH_8_33": value  <= 0.00321405893191695213;
            "FEATURE_THRESH_8_34": value  <= -0.00400232011452317238;
            "FEATURE_THRESH_8_35": value  <= 0.00741821294650435448;
            "FEATURE_THRESH_8_36": value  <= -0.00887645874172449112;
            "FEATURE_THRESH_8_37": value  <= 0.00273117399774491787;
            "FEATURE_THRESH_8_38": value  <= -0.00250823795795440674;
            "FEATURE_THRESH_8_39": value  <= -0.00805410742759704590;
            "FEATURE_THRESH_8_40": value  <= -0.00097938813269138336;
            "FEATURE_THRESH_8_41": value  <= -0.00587459094822406769;
            "FEATURE_THRESH_8_42": value  <= -0.00449367193505167961;
            "FEATURE_THRESH_8_43": value  <= -0.00543892290443181992;
            "FEATURE_THRESH_8_44": value  <= -0.00075094640487805009;
            "FEATURE_THRESH_8_45": value  <= 0.00001452880042052129;
            "FEATURE_THRESH_8_46": value  <= 0.04075806960463519701;
            "FEATURE_THRESH_8_47": value  <= 0.00665059313178062439;
            "FEATURE_THRESH_8_48": value  <= 0.00457593519240617752;
            "FEATURE_THRESH_8_49": value  <= 0.00652693118900060654;
            "FEATURE_THRESH_8_50": value  <= -0.01366037968546150033;
            "FEATURE_THRESH_8_51": value  <= 0.02735886909067630074;
            "FEATURE_THRESH_8_52": value  <= 0.00062197551596909761;
            "FEATURE_THRESH_8_53": value  <= -0.00330770807340741158;
            "FEATURE_THRESH_8_54": value  <= -0.01063110958784820037;
            "FEATURE_THRESH_8_55": value  <= 0.01944164931774140098;
            "FEATURE_THRESH_9_0": value  <= -0.00550521677359938622;
            "FEATURE_THRESH_9_1": value  <= 0.00195622793398797512;
            "FEATURE_THRESH_9_2": value  <= -0.00889247842133045197;
            "FEATURE_THRESH_9_3": value  <= 0.08363837748765949598;
            "FEATURE_THRESH_9_4": value  <= 0.00122822704724967480;
            "FEATURE_THRESH_9_5": value  <= 0.00576291698962450027;
            "FEATURE_THRESH_9_6": value  <= -0.00164174102246761322;
            "FEATURE_THRESH_9_7": value  <= 0.00341131491586565971;
            "FEATURE_THRESH_9_8": value  <= -0.01106932014226909983;
            "FEATURE_THRESH_9_9": value  <= 0.03486597165465350062;
            "FEATURE_THRESH_9_10": value  <= 0.00065701099811121821;
            "FEATURE_THRESH_9_11": value  <= -0.02433913014829160171;
            "FEATURE_THRESH_9_12": value  <= 0.00059435202274471521;
            "FEATURE_THRESH_9_13": value  <= 0.00229715090245008469;
            "FEATURE_THRESH_9_14": value  <= -0.00378018291667103767;
            "FEATURE_THRESH_9_15": value  <= -0.13420669734477999602;
            "FEATURE_THRESH_9_16": value  <= 0.00075224548345431685;
            "FEATURE_THRESH_9_17": value  <= -0.04054554179310800033;
            "FEATURE_THRESH_9_18": value  <= 0.00125729700084775686;
            "FEATURE_THRESH_9_19": value  <= -0.00742499483749270439;
            "FEATURE_THRESH_9_20": value  <= 0.00050908129196614027;
            "FEATURE_THRESH_9_21": value  <= -0.00128084502648562193;
            "FEATURE_THRESH_9_22": value  <= -0.00183488603215664625;
            "FEATURE_THRESH_9_23": value  <= 0.02748486958444119888;
            "FEATURE_THRESH_9_24": value  <= 0.00223724194802343845;
            "FEATURE_THRESH_9_25": value  <= -0.00886352919042110443;
            "FEATURE_THRESH_9_26": value  <= 0.00417539710178971291;
            "FEATURE_THRESH_9_27": value  <= -0.00170981895644217730;
            "FEATURE_THRESH_9_28": value  <= 0.00653285486623644829;
            "FEATURE_THRESH_9_29": value  <= -0.00953729078173637390;
            "FEATURE_THRESH_9_30": value  <= 0.02531098946928980048;
            "FEATURE_THRESH_9_31": value  <= 0.03646096959710119767;
            "FEATURE_THRESH_9_32": value  <= 0.02085432969033719844;
            "FEATURE_THRESH_9_33": value  <= -0.00087207747856155038;
            "FEATURE_THRESH_9_34": value  <= -0.00001522700040368363;
            "FEATURE_THRESH_9_35": value  <= -0.00084316509310156107;
            "FEATURE_THRESH_9_36": value  <= 0.00360378599725663662;
            "FEATURE_THRESH_9_37": value  <= -0.00680578919127583504;
            "FEATURE_THRESH_9_38": value  <= -0.04702166095376009852;
            "FEATURE_THRESH_9_39": value  <= -0.03695410862565039894;
            "FEATURE_THRESH_9_40": value  <= 0.00104394799564033747;
            "FEATURE_THRESH_9_41": value  <= -0.00021050689974799752;
            "FEATURE_THRESH_9_42": value  <= -0.08083158731460569901;
            "FEATURE_THRESH_9_43": value  <= -0.00036579059087671340;
            "FEATURE_THRESH_9_44": value  <= -0.00012545920617412776;
            "FEATURE_THRESH_9_45": value  <= -0.06878648698329929700;
            "FEATURE_THRESH_9_46": value  <= 0.01241578999906780070;
            "FEATURE_THRESH_9_47": value  <= -0.00471748178824782372;
            "FEATURE_THRESH_9_48": value  <= 0.03813685849308969672;
            "FEATURE_THRESH_9_49": value  <= -0.00281680491752922535;
            "FEATURE_THRESH_9_50": value  <= 0.00813036039471626282;
            "FEATURE_THRESH_9_51": value  <= 0.00600560195744037628;
            "FEATURE_THRESH_9_52": value  <= 0.01913931965827940160;
            "FEATURE_THRESH_9_53": value  <= 0.01644575968384739961;
            "FEATURE_THRESH_9_54": value  <= -0.03735689073801039956;
            "FEATURE_THRESH_9_55": value  <= -0.01972790062427520058;
            "FEATURE_THRESH_9_56": value  <= 0.00669725798070430756;
            "FEATURE_THRESH_9_57": value  <= 0.00074457528535276651;
            "FEATURE_THRESH_9_58": value  <= 0.00117906404193490744;
            "FEATURE_THRESH_9_59": value  <= 0.03498061001300809686;
            "FEATURE_THRESH_9_60": value  <= 0.00056859792675822973;
            "FEATURE_THRESH_9_61": value  <= -0.01134064979851250043;
            "FEATURE_THRESH_9_62": value  <= -0.00662281084805727005;
            "FEATURE_THRESH_9_63": value  <= -0.00801603309810161591;
            "FEATURE_THRESH_9_64": value  <= 0.00142068194691091776;
            "FEATURE_THRESH_9_65": value  <= -0.00278017111122608185;
            "FEATURE_THRESH_9_66": value  <= -0.00147475895937532187;
            "FEATURE_THRESH_9_67": value  <= -0.02383033931255339882;
            "FEATURE_THRESH_9_68": value  <= 0.00693697901442646980;
            "FEATURE_THRESH_9_69": value  <= 0.00828062556684017181;
            "FEATURE_THRESH_9_70": value  <= -0.01043950021266940031;
            "FEATURE_THRESH_10_0": value  <= 0.00720065878704190254;
            "FEATURE_THRESH_10_1": value  <= -0.00285935890860855579;
            "FEATURE_THRESH_10_2": value  <= 0.00068580528022721410;
            "FEATURE_THRESH_10_3": value  <= 0.00795801915228366852;
            "FEATURE_THRESH_10_4": value  <= -0.00121241505257785320;
            "FEATURE_THRESH_10_5": value  <= 0.00794261321425437927;
            "FEATURE_THRESH_10_6": value  <= 0.00246305903419852257;
            "FEATURE_THRESH_10_7": value  <= -0.00603965995833277702;
            "FEATURE_THRESH_10_8": value  <= -0.00129883398767560720;
            "FEATURE_THRESH_10_9": value  <= 0.00022299369447864592;
            "FEATURE_THRESH_10_10": value  <= 0.00146542803850024939;
            "FEATURE_THRESH_10_11": value  <= -0.00081210042117163539;
            "FEATURE_THRESH_10_12": value  <= -0.00138360203709453344;
            "FEATURE_THRESH_10_13": value  <= -0.02793644927442070006;
            "FEATURE_THRESH_10_14": value  <= -0.00046919551095925272;
            "FEATURE_THRESH_10_15": value  <= -0.00498296599835157394;
            "FEATURE_THRESH_10_16": value  <= 0.00188153097406029701;
            "FEATURE_THRESH_10_17": value  <= -0.01906755007803440094;
            "FEATURE_THRESH_10_18": value  <= -0.00469065597280859947;
            "FEATURE_THRESH_10_19": value  <= 0.00597771396860480309;
            "FEATURE_THRESH_10_20": value  <= -0.03330313041806220314;
            "FEATURE_THRESH_10_21": value  <= 0.09074410796165470472;
            "FEATURE_THRESH_10_22": value  <= 0.00093555898638442159;
            "FEATURE_THRESH_10_23": value  <= 0.01490165013819929989;
            "FEATURE_THRESH_10_24": value  <= 0.00061594118596985936;
            "FEATURE_THRESH_10_25": value  <= -0.05067098885774610345;
            "FEATURE_THRESH_10_26": value  <= 0.00068665749859064817;
            "FEATURE_THRESH_10_27": value  <= 0.00837124325335025787;
            "FEATURE_THRESH_10_28": value  <= -0.00129530695267021656;
            "FEATURE_THRESH_10_29": value  <= -0.04194168001413350194;
            "FEATURE_THRESH_10_30": value  <= -0.02352938055992129934;
            "FEATURE_THRESH_10_31": value  <= 0.04085744917392730019;
            "FEATURE_THRESH_10_32": value  <= -0.02540686912834640154;
            "FEATURE_THRESH_10_33": value  <= -0.00041415440500713885;
            "FEATURE_THRESH_10_34": value  <= 0.02182411961257460162;
            "FEATURE_THRESH_10_35": value  <= 0.01411403995007280004;
            "FEATURE_THRESH_10_36": value  <= 0.00006721459067193791;
            "FEATURE_THRESH_10_37": value  <= -0.00794176384806632996;
            "FEATURE_THRESH_10_38": value  <= -0.00721444096416234970;
            "FEATURE_THRESH_10_39": value  <= 0.00258173397742211819;
            "FEATURE_THRESH_10_40": value  <= 0.13409319519996640291;
            "FEATURE_THRESH_10_41": value  <= 0.00229627103544771671;
            "FEATURE_THRESH_10_42": value  <= -0.00215758499689400196;
            "FEATURE_THRESH_10_43": value  <= -0.00491961883381009102;
            "FEATURE_THRESH_10_44": value  <= 0.00162674696184694767;
            "FEATURE_THRESH_10_45": value  <= 0.00033413388882763684;
            "FEATURE_THRESH_10_46": value  <= -0.02669808082282540060;
            "FEATURE_THRESH_10_47": value  <= -0.03056187927722929867;
            "FEATURE_THRESH_10_48": value  <= 0.00285115488804876804;
            "FEATURE_THRESH_10_49": value  <= -0.03621147945523259942;
            "FEATURE_THRESH_10_50": value  <= -0.00241151894442737103;
            "FEATURE_THRESH_10_51": value  <= -0.00077253201743587852;
            "FEATURE_THRESH_10_52": value  <= 0.00029481729143299162;
            "FEATURE_THRESH_10_53": value  <= -0.00623345607891678810;
            "FEATURE_THRESH_10_54": value  <= -0.02627472952008250151;
            "FEATURE_THRESH_10_55": value  <= 0.00532122608274221420;
            "FEATURE_THRESH_10_56": value  <= -0.00411290582269430161;
            "FEATURE_THRESH_10_57": value  <= 0.00324578094296157360;
            "FEATURE_THRESH_10_58": value  <= -0.01635970920324330072;
            "FEATURE_THRESH_10_59": value  <= 0.00032166109303943813;
            "FEATURE_THRESH_10_60": value  <= 0.00064452440710738301;
            "FEATURE_THRESH_10_61": value  <= -0.00789097324013710022;
            "FEATURE_THRESH_10_62": value  <= 0.04833621159195899963;
            "FEATURE_THRESH_10_63": value  <= -0.00075178127735853195;
            "FEATURE_THRESH_10_64": value  <= -0.00249539106152951717;
            "FEATURE_THRESH_10_65": value  <= -0.00223850109614431858;
            "FEATURE_THRESH_10_66": value  <= -0.00179884303361177444;
            "FEATURE_THRESH_10_67": value  <= 0.00878609158098697662;
            "FEATURE_THRESH_10_68": value  <= 0.00367153808474540710;
            "FEATURE_THRESH_10_69": value  <= -0.03533644974231719971;
            "FEATURE_THRESH_10_70": value  <= -0.00069189240457490087;
            "FEATURE_THRESH_10_71": value  <= -0.00339461094699800014;
            "FEATURE_THRESH_10_72": value  <= 0.00098569283727556467;
            "FEATURE_THRESH_10_73": value  <= -0.05016310140490529840;
            "FEATURE_THRESH_10_74": value  <= -0.00223672599531710148;
            "FEATURE_THRESH_10_75": value  <= 0.00074326287722215056;
            "FEATURE_THRESH_10_76": value  <= -0.00093485182151198387;
            "FEATURE_THRESH_10_77": value  <= 0.01749793998897080163;
            "FEATURE_THRESH_10_78": value  <= -0.00152000004891306162;
            "FEATURE_THRESH_10_79": value  <= 0.00078003940870985389;
            "FEATURE_THRESH_11_0": value  <= -0.00999455526471138000;
            "FEATURE_THRESH_11_1": value  <= -0.00110852299258112907;
            "FEATURE_THRESH_11_2": value  <= 0.00103643804322928190;
            "FEATURE_THRESH_11_3": value  <= 0.00068211311008781195;
            "FEATURE_THRESH_11_4": value  <= -0.00068057340104132891;
            "FEATURE_THRESH_11_5": value  <= 0.00026068789884448051;
            "FEATURE_THRESH_11_6": value  <= 0.00051607372006401420;
            "FEATURE_THRESH_11_7": value  <= 0.00085007521556690335;
            "FEATURE_THRESH_11_8": value  <= -0.00186078296974301338;
            "FEATURE_THRESH_11_9": value  <= -0.00150339701212942600;
            "FEATURE_THRESH_11_10": value  <= 0.00234789098612964153;
            "FEATURE_THRESH_11_11": value  <= -0.00028880240279249847;
            "FEATURE_THRESH_11_12": value  <= 0.00894054770469665527;
            "FEATURE_THRESH_11_13": value  <= -0.01932773925364019915;
            "FEATURE_THRESH_11_14": value  <= -0.00020202060113660991;
            "FEATURE_THRESH_11_15": value  <= 0.00211790692992508411;
            "FEATURE_THRESH_11_16": value  <= -0.00177437602542340755;
            "FEATURE_THRESH_11_17": value  <= 0.00422344589605927467;
            "FEATURE_THRESH_11_18": value  <= -0.01437522005289790065;
            "FEATURE_THRESH_11_19": value  <= -0.01534918043762449960;
            "FEATURE_THRESH_11_20": value  <= 0.00001515227995696478;
            "FEATURE_THRESH_11_21": value  <= -0.00912939198315143585;
            "FEATURE_THRESH_11_22": value  <= 0.00225121597759425640;
            "FEATURE_THRESH_11_23": value  <= -0.00496969185769557953;
            "FEATURE_THRESH_11_24": value  <= -0.01282901037484410027;
            "FEATURE_THRESH_11_25": value  <= -0.00936600659042596817;
            "FEATURE_THRESH_11_26": value  <= 0.00324523192830383778;
            "FEATURE_THRESH_11_27": value  <= -0.01172356028109789935;
            "FEATURE_THRESH_11_28": value  <= 0.00002925794069597032;
            "FEATURE_THRESH_11_29": value  <= -0.00002224421950813849;
            "FEATURE_THRESH_11_30": value  <= 0.00508815096691250801;
            "FEATURE_THRESH_11_31": value  <= 0.02742967940866949950;
            "FEATURE_THRESH_11_32": value  <= -0.00641428679227828979;
            "FEATURE_THRESH_11_33": value  <= 0.00334799592383205891;
            "FEATURE_THRESH_11_34": value  <= -0.08263549208641049471;
            "FEATURE_THRESH_11_35": value  <= 0.00102617405354976654;
            "FEATURE_THRESH_11_36": value  <= -0.00163070904091000557;
            "FEATURE_THRESH_11_37": value  <= 0.00245466805063188076;
            "FEATURE_THRESH_11_38": value  <= -0.00099476519972085953;
            "FEATURE_THRESH_11_39": value  <= 0.01540919020771979939;
            "FEATURE_THRESH_11_40": value  <= 0.00117844005580991507;
            "FEATURE_THRESH_11_41": value  <= -0.02770191989839080118;
            "FEATURE_THRESH_11_42": value  <= -0.02950539998710159997;
            "FEATURE_THRESH_11_43": value  <= 0.00045159430010244250;
            "FEATURE_THRESH_11_44": value  <= 0.00717726396396756172;
            "FEATURE_THRESH_11_45": value  <= -0.07418204843997959486;
            "FEATURE_THRESH_11_46": value  <= -0.01725416071712970040;
            "FEATURE_THRESH_11_47": value  <= 0.01485155988484620007;
            "FEATURE_THRESH_11_48": value  <= 0.01000200025737289951;
            "FEATURE_THRESH_11_49": value  <= 0.00201381207443773746;
            "FEATURE_THRESH_11_50": value  <= 0.00151354703120887280;
            "FEATURE_THRESH_11_51": value  <= 0.00313814310356974602;
            "FEATURE_THRESH_11_52": value  <= -0.00514504406601190567;
            "FEATURE_THRESH_11_53": value  <= -0.00447367085143923759;
            "FEATURE_THRESH_11_54": value  <= 0.00196284707635641098;
            "FEATURE_THRESH_11_55": value  <= 0.00542604504153132439;
            "FEATURE_THRESH_11_56": value  <= 0.00049611460417509079;
            "FEATURE_THRESH_11_57": value  <= 0.00937287881970405579;
            "FEATURE_THRESH_11_58": value  <= 0.00060500897234305739;
            "FEATURE_THRESH_11_59": value  <= 0.00056792551185935736;
            "FEATURE_THRESH_11_60": value  <= 0.02464433945715429827;
            "FEATURE_THRESH_11_61": value  <= -0.01029045041650530033;
            "FEATURE_THRESH_11_62": value  <= 0.00206294190138578415;
            "FEATURE_THRESH_11_63": value  <= -0.00505194813013076782;
            "FEATURE_THRESH_11_64": value  <= -0.00576926209032535553;
            "FEATURE_THRESH_11_65": value  <= -0.00045789941214025021;
            "FEATURE_THRESH_11_66": value  <= -0.00075918837683275342;
            "FEATURE_THRESH_11_67": value  <= -0.00177372596226632595;
            "FEATURE_THRESH_11_68": value  <= -0.00856104679405689240;
            "FEATURE_THRESH_11_69": value  <= 0.00172772700898349285;
            "FEATURE_THRESH_11_70": value  <= -0.02819960936903950083;
            "FEATURE_THRESH_11_71": value  <= -0.00177811097819358110;
            "FEATURE_THRESH_11_72": value  <= 0.00033177141449414194;
            "FEATURE_THRESH_11_73": value  <= 0.00263853999786078930;
            "FEATURE_THRESH_11_74": value  <= -0.00211830693297088146;
            "FEATURE_THRESH_11_75": value  <= -0.01477328967303040072;
            "FEATURE_THRESH_11_76": value  <= -0.01681544072926039954;
            "FEATURE_THRESH_11_77": value  <= -0.00633701402693986893;
            "FEATURE_THRESH_11_78": value  <= -0.00004456004899111577;
            "FEATURE_THRESH_11_79": value  <= -0.00102406204678118229;
            "FEATURE_THRESH_11_80": value  <= -0.00231616897508502007;
            "FEATURE_THRESH_11_81": value  <= 0.53217571973800659180;
            "FEATURE_THRESH_11_82": value  <= -0.16643050312995910645;
            "FEATURE_THRESH_11_83": value  <= 0.11253529787063600021;
            "FEATURE_THRESH_11_84": value  <= 0.00930468644946813583;
            "FEATURE_THRESH_11_85": value  <= -0.00462550995871424675;
            "FEATURE_THRESH_11_86": value  <= -0.11116469651460650359;
            "FEATURE_THRESH_11_87": value  <= -0.01088843960314989957;
            "FEATURE_THRESH_11_88": value  <= 0.00585643015801906586;
            "FEATURE_THRESH_11_89": value  <= 0.05485438928008080223;
            "FEATURE_THRESH_11_90": value  <= -0.01119733974337580075;
            "FEATURE_THRESH_11_91": value  <= 0.00440690713003277779;
            "FEATURE_THRESH_11_92": value  <= -0.06366529315710070525;
            "FEATURE_THRESH_11_93": value  <= -0.00980814918875694275;
            "FEATURE_THRESH_11_94": value  <= -0.00217170990072190762;
            "FEATURE_THRESH_11_95": value  <= -0.01331552024930720071;
            "FEATURE_THRESH_11_96": value  <= 0.00254420796409249306;
            "FEATURE_THRESH_11_97": value  <= 0.01203783974051480035;
            "FEATURE_THRESH_11_98": value  <= -0.02070105075836179906;
            "FEATURE_THRESH_11_99": value  <= 0.02760827913880349940;
            "FEATURE_THRESH_11_100": value  <= 0.00123706203885376453;
            "FEATURE_THRESH_11_101": value  <= -0.03766933828592299721;
            "FEATURE_THRESH_11_102": value  <= -0.00180572597309947014;
            "FEATURE_THRESH_12_0": value  <= 0.00442990288138389587;
            "FEATURE_THRESH_12_1": value  <= -0.00238133198581635952;
            "FEATURE_THRESH_12_2": value  <= 0.00229157111607491970;
            "FEATURE_THRESH_12_3": value  <= 0.00099457940086722374;
            "FEATURE_THRESH_12_4": value  <= 0.00077164667891338468;
            "FEATURE_THRESH_12_5": value  <= -0.00113864103332161903;
            "FEATURE_THRESH_12_6": value  <= -0.00016403039626311511;
            "FEATURE_THRESH_12_7": value  <= 0.00002979352939291858;
            "FEATURE_THRESH_12_8": value  <= 0.00857749022543430328;
            "FEATURE_THRESH_12_9": value  <= -0.00026032689493149519;
            "FEATURE_THRESH_12_10": value  <= -0.00614046305418014526;
            "FEATURE_THRESH_12_11": value  <= -0.02308695018291469919;
            "FEATURE_THRESH_12_12": value  <= -0.01424365025013690084;
            "FEATURE_THRESH_12_13": value  <= 0.01948712952435020102;
            "FEATURE_THRESH_12_14": value  <= -0.00096681108698248863;
            "FEATURE_THRESH_12_15": value  <= 0.00314747099764645100;
            "FEATURE_THRESH_12_16": value  <= -0.00018026070029009134;
            "FEATURE_THRESH_12_17": value  <= -0.00602662609890103340;
            "FEATURE_THRESH_12_18": value  <= 0.00044462960795499384;
            "FEATURE_THRESH_12_19": value  <= 0.00226097600534558296;
            "FEATURE_THRESH_12_20": value  <= 0.05113305896520609767;
            "FEATURE_THRESH_12_21": value  <= -0.01778630912303920050;
            "FEATURE_THRESH_12_22": value  <= -0.00496796285733580589;
            "FEATURE_THRESH_12_23": value  <= 0.00206676893867552280;
            "FEATURE_THRESH_12_24": value  <= 0.00744137680158019066;
            "FEATURE_THRESH_12_25": value  <= -0.00362772797234356403;
            "FEATURE_THRESH_12_26": value  <= -0.00535307591781020164;
            "FEATURE_THRESH_12_27": value  <= 0.14530919492244720459;
            "FEATURE_THRESH_12_28": value  <= 0.00243944907560944557;
            "FEATURE_THRESH_12_29": value  <= -0.00312833907082676888;
            "FEATURE_THRESH_12_30": value  <= 0.00179402600042521954;
            "FEATURE_THRESH_12_31": value  <= 0.03625382110476489672;
            "FEATURE_THRESH_12_32": value  <= -0.00517467223107814789;
            "FEATURE_THRESH_12_33": value  <= 0.00065383297624066472;
            "FEATURE_THRESH_12_34": value  <= -0.02648022957146169837;
            "FEATURE_THRESH_12_35": value  <= -0.00304406601935625076;
            "FEATURE_THRESH_12_36": value  <= 0.00369935203343629837;
            "FEATURE_THRESH_12_37": value  <= -0.00036762931267730892;
            "FEATURE_THRESH_12_38": value  <= -0.04138226062059399690;
            "FEATURE_THRESH_12_39": value  <= -0.00105327297933399677;
            "FEATURE_THRESH_12_40": value  <= -0.00216486002318561077;
            "FEATURE_THRESH_12_41": value  <= -0.00056747748749330640;
            "FEATURE_THRESH_12_42": value  <= 0.17375840246677398682;
            "FEATURE_THRESH_12_43": value  <= -0.00290496996603906155;
            "FEATURE_THRESH_12_44": value  <= 0.00122995395213365555;
            "FEATURE_THRESH_12_45": value  <= -0.00054329237900674343;
            "FEATURE_THRESH_12_46": value  <= -0.00832972582429647446;
            "FEATURE_THRESH_12_47": value  <= -0.00010417630255687982;
            "FEATURE_THRESH_12_48": value  <= 0.03120470046997069966;
            "FEATURE_THRESH_12_49": value  <= 0.00789435021579265594;
            "FEATURE_THRESH_12_50": value  <= -0.00436453102156519890;
            "FEATURE_THRESH_12_51": value  <= 0.00767930597066879272;
            "FEATURE_THRESH_12_52": value  <= -0.02543113939464090173;
            "FEATURE_THRESH_12_53": value  <= 0.00082000601105391979;
            "FEATURE_THRESH_12_54": value  <= 0.00292846001684665680;
            "FEATURE_THRESH_12_55": value  <= 0.00004525647091213614;
            "FEATURE_THRESH_12_56": value  <= 0.00131583097390830517;
            "FEATURE_THRESH_12_57": value  <= 0.00158703897614032030;
            "FEATURE_THRESH_12_58": value  <= -0.02153966017067429975;
            "FEATURE_THRESH_12_59": value  <= 0.01433448027819399923;
            "FEATURE_THRESH_12_60": value  <= -0.00838813837617635727;
            "FEATURE_THRESH_12_61": value  <= 0.00919068418443202972;
            "FEATURE_THRESH_12_62": value  <= -0.00584530597552657127;
            "FEATURE_THRESH_12_63": value  <= -0.05470779910683629815;
            "FEATURE_THRESH_12_64": value  <= 0.00911427754908800125;
            "FEATURE_THRESH_12_65": value  <= -0.01557500008493659972;
            "FEATURE_THRESH_12_66": value  <= -0.00012050600344082341;
            "FEATURE_THRESH_12_67": value  <= 0.00122739700600504875;
            "FEATURE_THRESH_12_68": value  <= -0.00121866003610193729;
            "FEATURE_THRESH_12_69": value  <= -0.00332566490396857262;
            "FEATURE_THRESH_12_70": value  <= -0.01328830979764459956;
            "FEATURE_THRESH_12_71": value  <= -0.00338397710584104061;
            "FEATURE_THRESH_12_72": value  <= -0.21954220533370968904;
            "FEATURE_THRESH_12_73": value  <= 0.00491117080673575401;
            "FEATURE_THRESH_12_74": value  <= -0.00018744950648397207;
            "FEATURE_THRESH_12_75": value  <= -0.00521786417812108994;
            "FEATURE_THRESH_12_76": value  <= -0.00111115199979394674;
            "FEATURE_THRESH_12_77": value  <= 0.00440364005044102669;
            "FEATURE_THRESH_12_78": value  <= 0.12299499660730360551;
            "FEATURE_THRESH_12_79": value  <= -0.01231351029127840044;
            "FEATURE_THRESH_12_80": value  <= 0.00414710398763418198;
            "FEATURE_THRESH_12_81": value  <= -0.00355026498436927795;
            "FEATURE_THRESH_12_82": value  <= -0.01922426931560039867;
            "FEATURE_THRESH_12_83": value  <= 0.00143950595520436764;
            "FEATURE_THRESH_12_84": value  <= -0.00677519990131258965;
            "FEATURE_THRESH_12_85": value  <= 0.00701196305453777313;
            "FEATURE_THRESH_12_86": value  <= 0.00540146511048078537;
            "FEATURE_THRESH_12_87": value  <= 0.00090274988906458020;
            "FEATURE_THRESH_12_88": value  <= 0.01147445011883970085;
            "FEATURE_THRESH_12_89": value  <= -0.00670234300196170807;
            "FEATURE_THRESH_12_90": value  <= -0.00204629590734839439;
            "FEATURE_THRESH_12_91": value  <= -0.00999515689909458160;
            "FEATURE_THRESH_12_92": value  <= -0.03570070862770079873;
            "FEATURE_THRESH_12_93": value  <= 0.00045584561303257942;
            "FEATURE_THRESH_12_94": value  <= -0.05426060035824779859;
            "FEATURE_THRESH_12_95": value  <= 0.00606004614382982254;
            "FEATURE_THRESH_12_96": value  <= -0.00647918321192264557;
            "FEATURE_THRESH_12_97": value  <= -0.00149394699838012457;
            "FEATURE_THRESH_12_98": value  <= 0.00001461053034290672;
            "FEATURE_THRESH_12_99": value  <= -0.00723219383507966995;
            "FEATURE_THRESH_12_100": value  <= -0.00406458182260394096;
            "FEATURE_THRESH_12_101": value  <= 0.03046308085322380066;
            "FEATURE_THRESH_12_102": value  <= -0.00805449113249778748;
            "FEATURE_THRESH_12_103": value  <= 0.03950513899326320300;
            "FEATURE_THRESH_12_104": value  <= 0.00845302082598209381;
            "FEATURE_THRESH_12_105": value  <= -0.00116881204303354025;
            "FEATURE_THRESH_12_106": value  <= 0.00280706700868904591;
            "FEATURE_THRESH_12_107": value  <= 0.00047365209320560098;
            "FEATURE_THRESH_12_108": value  <= 0.01174108032137160043;
            "FEATURE_THRESH_12_109": value  <= 0.00318332388997077942;
            "FEATURE_THRESH_12_110": value  <= 0.00070241501089185476;
            "FEATURE_THRESH_13_0": value  <= 0.01705992966890339940;
            "FEATURE_THRESH_13_1": value  <= 0.02184084057807919935;
            "FEATURE_THRESH_13_2": value  <= 0.00024520049919374287;
            "FEATURE_THRESH_13_3": value  <= 0.00832726061344146729;
            "FEATURE_THRESH_13_4": value  <= 0.00057148298947140574;
            "FEATURE_THRESH_13_5": value  <= 0.00067373987985774875;
            "FEATURE_THRESH_13_6": value  <= 0.00003468159047770314;
            "FEATURE_THRESH_13_7": value  <= -0.00585633981972932816;
            "FEATURE_THRESH_13_8": value  <= 0.00851022731512784958;
            "FEATURE_THRESH_13_9": value  <= -0.06981720775365829468;
            "FEATURE_THRESH_13_10": value  <= -0.00086113670840859413;
            "FEATURE_THRESH_13_11": value  <= 0.00097149249631911516;
            "FEATURE_THRESH_13_12": value  <= -0.00001472749045206001;
            "FEATURE_THRESH_13_13": value  <= 0.04842029139399529891;
            "FEATURE_THRESH_13_14": value  <= 0.00132571405265480280;
            "FEATURE_THRESH_13_15": value  <= 0.00001492214960308047;
            "FEATURE_THRESH_13_16": value  <= -0.00271733989939093590;
            "FEATURE_THRESH_13_17": value  <= 0.00292195007205009460;
            "FEATURE_THRESH_13_18": value  <= -0.00198049889877438545;
            "FEATURE_THRESH_13_19": value  <= -0.00400121090933680534;
            "FEATURE_THRESH_13_20": value  <= -0.00434919912368059158;
            "FEATURE_THRESH_13_21": value  <= 0.00134908896870911121;
            "FEATURE_THRESH_13_22": value  <= 0.01859707012772560120;
            "FEATURE_THRESH_13_23": value  <= -0.00185623799916356802;
            "FEATURE_THRESH_13_24": value  <= 0.00229404307901859283;
            "FEATURE_THRESH_13_25": value  <= 0.00029982850537635386;
            "FEATURE_THRESH_13_26": value  <= 0.00354554597288370132;
            "FEATURE_THRESH_13_27": value  <= 0.00961047224700450897;
            "FEATURE_THRESH_13_28": value  <= -0.00627832207828760147;
            "FEATURE_THRESH_13_29": value  <= 0.00345984799787402153;
            "FEATURE_THRESH_13_30": value  <= -0.00131120195146650076;
            "FEATURE_THRESH_13_31": value  <= 0.00268761790357530117;
            "FEATURE_THRESH_13_32": value  <= 0.00391181698068976402;
            "FEATURE_THRESH_13_33": value  <= -0.01420645043253900008;
            "FEATURE_THRESH_13_34": value  <= 0.00071705528534948826;
            "FEATURE_THRESH_13_35": value  <= 0.00166350195650011301;
            "FEATURE_THRESH_13_36": value  <= 0.00336861889809370041;
            "FEATURE_THRESH_13_37": value  <= 0.01279953029006719936;
            "FEATURE_THRESH_13_38": value  <= 0.00339012010954320431;
            "FEATURE_THRESH_13_39": value  <= 0.00470707798376679420;
            "FEATURE_THRESH_13_40": value  <= 0.00148193398490548134;
            "FEATURE_THRESH_13_41": value  <= -0.00699957599863409996;
            "FEATURE_THRESH_13_42": value  <= 0.01593901030719279896;
            "FEATURE_THRESH_13_43": value  <= 0.00763773499056696892;
            "FEATURE_THRESH_13_44": value  <= 0.00673340400680899620;
            "FEATURE_THRESH_13_45": value  <= -0.01285880990326400061;
            "FEATURE_THRESH_13_46": value  <= -0.00062270800117403269;
            "FEATURE_THRESH_13_47": value  <= -0.00052651681471616030;
            "FEATURE_THRESH_13_48": value  <= 0.01107509993016719992;
            "FEATURE_THRESH_13_49": value  <= -0.03672825172543529859;
            "FEATURE_THRESH_13_50": value  <= -0.00028207109426148236;
            "FEATURE_THRESH_13_51": value  <= -0.00274896901100873947;
            "FEATURE_THRESH_13_52": value  <= 0.01004751957952980043;
            "FEATURE_THRESH_13_53": value  <= -0.00814978405833244324;
            "FEATURE_THRESH_13_54": value  <= -0.00688338885083794594;
            "FEATURE_THRESH_13_55": value  <= -0.00001403936039423570;
            "FEATURE_THRESH_13_56": value  <= 0.00154984195251017809;
            "FEATURE_THRESH_13_57": value  <= -0.00678414991125464439;
            "FEATURE_THRESH_13_58": value  <= 0.00021705629478674382;
            "FEATURE_THRESH_13_59": value  <= 0.00031198898795992136;
            "FEATURE_THRESH_13_60": value  <= 0.00545075302943587303;
            "FEATURE_THRESH_13_61": value  <= -0.00025818689027801156;
            "FEATURE_THRESH_13_62": value  <= -0.01744253933429720099;
            "FEATURE_THRESH_13_63": value  <= -0.04534352943301200173;
            "FEATURE_THRESH_13_64": value  <= 0.00191906897816807032;
            "FEATURE_THRESH_13_65": value  <= -0.00601778691634535789;
            "FEATURE_THRESH_13_66": value  <= -0.00407207384705543518;
            "FEATURE_THRESH_13_67": value  <= 0.00039855059003457427;
            "FEATURE_THRESH_13_68": value  <= -0.00654185703024268150;
            "FEATURE_THRESH_13_69": value  <= 0.00348450895398855209;
            "FEATURE_THRESH_13_70": value  <= -0.01369678042829040009;
            "FEATURE_THRESH_13_71": value  <= -0.01734714023768900090;
            "FEATURE_THRESH_13_72": value  <= -0.00408854288980364799;
            "FEATURE_THRESH_13_73": value  <= -0.00946879014372825623;
            "FEATURE_THRESH_13_74": value  <= 0.00170848402194678783;
            "FEATURE_THRESH_13_75": value  <= 0.00948090944439172745;
            "FEATURE_THRESH_13_76": value  <= -0.00473896507173776627;
            "FEATURE_THRESH_13_77": value  <= 0.00657610502094030380;
            "FEATURE_THRESH_13_78": value  <= -0.00216905493289232254;
            "FEATURE_THRESH_13_79": value  <= 0.01466017030179500059;
            "FEATURE_THRESH_13_80": value  <= 0.00017231999663636088;
            "FEATURE_THRESH_13_81": value  <= -0.02180376090109350032;
            "FEATURE_THRESH_13_82": value  <= -0.09473610669374470106;
            "FEATURE_THRESH_13_83": value  <= 0.00558255519717931747;
            "FEATURE_THRESH_13_84": value  <= 0.00195170904044061899;
            "FEATURE_THRESH_13_85": value  <= 0.01214990019798280023;
            "FEATURE_THRESH_13_86": value  <= -0.00751696201041340828;
            "FEATURE_THRESH_13_87": value  <= -0.07166790962219239669;
            "FEATURE_THRESH_13_88": value  <= -0.08829241991043089433;
            "FEATURE_THRESH_13_89": value  <= 0.03106307983398439929;
            "FEATURE_THRESH_13_90": value  <= 0.04662184044718740289;
            "FEATURE_THRESH_13_91": value  <= -0.01218948978930710011;
            "FEATURE_THRESH_13_92": value  <= 0.01301611028611660004;
            "FEATURE_THRESH_13_93": value  <= -0.00349528994411230087;
            "FEATURE_THRESH_13_94": value  <= -0.00004401503974804655;
            "FEATURE_THRESH_13_95": value  <= -0.10966490209102630615;
            "FEATURE_THRESH_13_96": value  <= -0.00090279558207839727;
            "FEATURE_THRESH_13_97": value  <= 0.00071126641705632210;
            "FEATURE_THRESH_13_98": value  <= -0.00312502798624336720;
            "FEATURE_THRESH_13_99": value  <= 0.00241446797735989094;
            "FEATURE_THRESH_13_100": value  <= 0.00044391240226104856;
            "FEATURE_THRESH_13_101": value  <= -0.00022611189342569560;
            "FEATURE_THRESH_14_0": value  <= -0.04690128937363619716;
            "FEATURE_THRESH_14_1": value  <= -0.00145683495793491602;
            "FEATURE_THRESH_14_2": value  <= 0.00555983697995543480;
            "FEATURE_THRESH_14_3": value  <= 0.00073170487303286791;
            "FEATURE_THRESH_14_4": value  <= 0.00133180094417184591;
            "FEATURE_THRESH_14_5": value  <= 0.00024347059661522508;
            "FEATURE_THRESH_14_6": value  <= -0.00305124698206782341;
            "FEATURE_THRESH_14_7": value  <= -0.00068657199153676629;
            "FEATURE_THRESH_14_8": value  <= 0.00146682001650333405;
            "FEATURE_THRESH_14_9": value  <= 0.00032021870720200241;
            "FEATURE_THRESH_14_10": value  <= 0.00074122188379988074;
            "FEATURE_THRESH_14_11": value  <= 0.00383302988484501839;
            "FEATURE_THRESH_14_12": value  <= -0.01545643992722029944;
            "FEATURE_THRESH_14_13": value  <= 0.00267967791296541691;
            "FEATURE_THRESH_14_14": value  <= 0.00282965693622827530;
            "FEATURE_THRESH_14_15": value  <= -0.00394442491233348846;
            "FEATURE_THRESH_14_16": value  <= 0.00271795596927404404;
            "FEATURE_THRESH_14_17": value  <= 0.00590776279568672180;
            "FEATURE_THRESH_14_18": value  <= -0.00422403495758771896;
            "FEATURE_THRESH_14_19": value  <= 0.00407258886843919754;
            "FEATURE_THRESH_14_20": value  <= 0.01014953013509510039;
            "FEATURE_THRESH_14_21": value  <= -0.00018864999583456665;
            "FEATURE_THRESH_14_22": value  <= -0.00488643581047654152;
            "FEATURE_THRESH_14_23": value  <= 0.02615847997367379968;
            "FEATURE_THRESH_14_24": value  <= 0.00048560759751126170;
            "FEATURE_THRESH_14_25": value  <= 0.01126870978623630004;
            "FEATURE_THRESH_14_26": value  <= -0.00281146191991865635;
            "FEATURE_THRESH_14_27": value  <= -0.00561127299442887306;
            "FEATURE_THRESH_14_28": value  <= 0.00856800936162471771;
            "FEATURE_THRESH_14_29": value  <= -0.00038172779022715986;
            "FEATURE_THRESH_14_30": value  <= -0.00017680290329735726;
            "FEATURE_THRESH_14_31": value  <= 0.00651125377044081688;
            "FEATURE_THRESH_14_32": value  <= -0.00006594868318643421;
            "FEATURE_THRESH_14_33": value  <= 0.00699390517547726631;
            "FEATURE_THRESH_14_34": value  <= -0.00467444397509098053;
            "FEATURE_THRESH_14_35": value  <= 0.01158985029906029959;
            "FEATURE_THRESH_14_36": value  <= 0.01300784014165400071;
            "FEATURE_THRESH_14_37": value  <= -0.00110085797496140003;
            "FEATURE_THRESH_14_38": value  <= 0.00060472649056464434;
            "FEATURE_THRESH_14_39": value  <= -0.01449484005570409947;
            "FEATURE_THRESH_14_40": value  <= -0.00530569488182663918;
            "FEATURE_THRESH_14_41": value  <= -0.00081829127157106996;
            "FEATURE_THRESH_14_42": value  <= -0.01907752081751819956;
            "FEATURE_THRESH_14_43": value  <= 0.00035549470339901745;
            "FEATURE_THRESH_14_44": value  <= 0.00196797307580709457;
            "FEATURE_THRESH_14_45": value  <= 0.00691891415044665337;
            "FEATURE_THRESH_14_46": value  <= 0.00298727792687714100;
            "FEATURE_THRESH_14_47": value  <= -0.00622646184638142586;
            "FEATURE_THRESH_14_48": value  <= 0.01335330028086900017;
            "FEATURE_THRESH_14_49": value  <= 0.03350523859262469900;
            "FEATURE_THRESH_14_50": value  <= -0.00252944603562355042;
            "FEATURE_THRESH_14_51": value  <= -0.00128016294911503792;
            "FEATURE_THRESH_14_52": value  <= 0.00706873880699276924;
            "FEATURE_THRESH_14_53": value  <= 0.00096880499040707946;
            "FEATURE_THRESH_14_54": value  <= 0.00396476592868566513;
            "FEATURE_THRESH_14_55": value  <= -0.02205773070454599902;
            "FEATURE_THRESH_14_56": value  <= -0.00066906312713399529;
            "FEATURE_THRESH_14_57": value  <= -0.00067009328631684184;
            "FEATURE_THRESH_14_58": value  <= 0.00074284552829340100;
            "FEATURE_THRESH_14_59": value  <= 0.00222278106957674026;
            "FEATURE_THRESH_14_60": value  <= -0.00541305216029286385;
            "FEATURE_THRESH_14_61": value  <= -0.00001452004016755382;
            "FEATURE_THRESH_14_62": value  <= 0.00023369169502984732;
            "FEATURE_THRESH_14_63": value  <= 0.00428945478051900864;
            "FEATURE_THRESH_14_64": value  <= 0.00591031508520245552;
            "FEATURE_THRESH_14_65": value  <= 0.01290053967386479983;
            "FEATURE_THRESH_14_66": value  <= 0.00469829794019460678;
            "FEATURE_THRESH_14_67": value  <= 0.01043985970318320015;
            "FEATURE_THRESH_14_68": value  <= 0.00304431910626590252;
            "FEATURE_THRESH_14_69": value  <= -0.00061593751888722181;
            "FEATURE_THRESH_14_70": value  <= -0.00342471594922244549;
            "FEATURE_THRESH_14_71": value  <= -0.00935385655611753464;
            "FEATURE_THRESH_14_72": value  <= 0.05233899876475330004;
            "FEATURE_THRESH_14_73": value  <= 0.00357656204141676426;
            "FEATURE_THRESH_14_74": value  <= 0.00071555317845195532;
            "FEATURE_THRESH_14_75": value  <= -0.01051667984575030065;
            "FEATURE_THRESH_14_76": value  <= 0.00773479277268052101;
            "FEATURE_THRESH_14_77": value  <= -0.00432267785072326660;
            "FEATURE_THRESH_14_78": value  <= -0.00255343993194401264;
            "FEATURE_THRESH_14_79": value  <= 0.00010268510231981054;
            "FEATURE_THRESH_14_80": value  <= 0.00000713951885700226;
            "FEATURE_THRESH_14_81": value  <= -0.00167119898833334446;
            "FEATURE_THRESH_14_82": value  <= 0.00492604495957493782;
            "FEATURE_THRESH_14_83": value  <= 0.00439087022095918655;
            "FEATURE_THRESH_14_84": value  <= -0.01779362931847569898;
            "FEATURE_THRESH_14_85": value  <= 0.00204696692526340485;
            "FEATURE_THRESH_14_86": value  <= 0.02989148907363409907;
            "FEATURE_THRESH_14_87": value  <= 0.00154949002899229527;
            "FEATURE_THRESH_14_88": value  <= 0.00149569695349782705;
            "FEATURE_THRESH_14_89": value  <= 0.00095885928021743894;
            "FEATURE_THRESH_14_90": value  <= 0.00049643701640889049;
            "FEATURE_THRESH_14_91": value  <= -0.00272808107547461987;
            "FEATURE_THRESH_14_92": value  <= 0.00230264803394675255;
            "FEATURE_THRESH_14_93": value  <= 0.25151631236076360532;
            "FEATURE_THRESH_14_94": value  <= -0.00463280221447348595;
            "FEATURE_THRESH_14_95": value  <= -0.04043449088931080210;
            "FEATURE_THRESH_14_96": value  <= 0.00001497222001489718;
            "FEATURE_THRESH_14_97": value  <= -0.00024050309730228037;
            "FEATURE_THRESH_14_98": value  <= 0.02365783974528309908;
            "FEATURE_THRESH_14_99": value  <= -0.00814491044729948044;
            "FEATURE_THRESH_14_100": value  <= -0.00369921303354203701;
            "FEATURE_THRESH_14_101": value  <= -0.00677186017856001854;
            "FEATURE_THRESH_14_102": value  <= 0.00426695309579372406;
            "FEATURE_THRESH_14_103": value  <= 0.00177919899579137564;
            "FEATURE_THRESH_14_104": value  <= 0.00167747703380882740;
            "FEATURE_THRESH_14_105": value  <= 0.00117326295003294945;
            "FEATURE_THRESH_14_106": value  <= 0.00086998171173036098;
            "FEATURE_THRESH_14_107": value  <= 0.00076378340600058436;
            "FEATURE_THRESH_14_108": value  <= 0.00015684569370932877;
            "FEATURE_THRESH_14_109": value  <= -0.02151137031614780079;
            "FEATURE_THRESH_14_110": value  <= 0.00013081369979772717;
            "FEATURE_THRESH_14_111": value  <= 0.02199204079806800147;
            "FEATURE_THRESH_14_112": value  <= -0.00080136500764638186;
            "FEATURE_THRESH_14_113": value  <= -0.00827360991388559341;
            "FEATURE_THRESH_14_114": value  <= 0.00368317891843616962;
            "FEATURE_THRESH_14_115": value  <= -0.00795256812125444412;
            "FEATURE_THRESH_14_116": value  <= 0.00153822998981922865;
            "FEATURE_THRESH_14_117": value  <= -0.01404353044927120035;
            "FEATURE_THRESH_14_118": value  <= 0.00143158901482820511;
            "FEATURE_THRESH_14_119": value  <= -0.03401422873139380021;
            "FEATURE_THRESH_14_120": value  <= -0.01202729996293780065;
            "FEATURE_THRESH_14_121": value  <= 0.13316619396209719572;
            "FEATURE_THRESH_14_122": value  <= -0.00152219494339078665;
            "FEATURE_THRESH_14_123": value  <= -0.00093929271679371595;
            "FEATURE_THRESH_14_124": value  <= 0.02771973982453350069;
            "FEATURE_THRESH_14_125": value  <= 0.00310301501303911209;
            "FEATURE_THRESH_14_126": value  <= 0.07786121964454649491;
            "FEATURE_THRESH_14_127": value  <= -0.01585493981838230135;
            "FEATURE_THRESH_14_128": value  <= -0.00497253006324172020;
            "FEATURE_THRESH_14_129": value  <= -0.00097676506265997887;
            "FEATURE_THRESH_14_130": value  <= -0.00246477103792130947;
            "FEATURE_THRESH_14_131": value  <= -0.00679377000778913498;
            "FEATURE_THRESH_14_132": value  <= 0.03260802105069159768;
            "FEATURE_THRESH_14_133": value  <= -0.00058514421107247472;
            "FEATURE_THRESH_14_134": value  <= -0.02963260002434249876;
            "FEATURE_THRESH_15_0": value  <= 0.04655085131525989878;
            "FEATURE_THRESH_15_1": value  <= 0.00795371271669864655;
            "FEATURE_THRESH_15_2": value  <= 0.00068221561377868056;
            "FEATURE_THRESH_15_3": value  <= -0.00019348249770700932;
            "FEATURE_THRESH_15_4": value  <= -0.00026710508973337710;
            "FEATURE_THRESH_15_5": value  <= 0.00278180604800581932;
            "FEATURE_THRESH_15_6": value  <= -0.00046779078547842801;
            "FEATURE_THRESH_15_7": value  <= -0.00003033516077266541;
            "FEATURE_THRESH_15_8": value  <= 0.00078038009814918041;
            "FEATURE_THRESH_15_9": value  <= -0.00425538513809442520;
            "FEATURE_THRESH_15_10": value  <= -0.00024735610350035131;
            "FEATURE_THRESH_15_11": value  <= -0.00014724259381182492;
            "FEATURE_THRESH_15_12": value  <= 0.00118647702038288116;
            "FEATURE_THRESH_15_13": value  <= 0.00239365804009139538;
            "FEATURE_THRESH_15_14": value  <= -0.00153905397746711969;
            "FEATURE_THRESH_15_15": value  <= -0.00719687901437282562;
            "FEATURE_THRESH_15_16": value  <= -0.00041499789222143590;
            "FEATURE_THRESH_15_17": value  <= 0.00443598302081227303;
            "FEATURE_THRESH_15_18": value  <= 0.00266062002629041672;
            "FEATURE_THRESH_15_19": value  <= -0.00152872002217918634;
            "FEATURE_THRESH_15_20": value  <= -0.00473972503095865250;
            "FEATURE_THRESH_15_21": value  <= -0.01482912991195920079;
            "FEATURE_THRESH_15_22": value  <= 0.00092275557108223438;
            "FEATURE_THRESH_15_23": value  <= 0.08352980762720109420;
            "FEATURE_THRESH_15_24": value  <= -0.00075633148662745953;
            "FEATURE_THRESH_15_25": value  <= 0.00984038598835468292;
            "FEATURE_THRESH_15_26": value  <= -0.00159538304433226585;
            "FEATURE_THRESH_15_27": value  <= 0.00003476602068985812;
            "FEATURE_THRESH_15_28": value  <= 0.02986291050910950054;
            "FEATURE_THRESH_15_29": value  <= 0.01132559031248090049;
            "FEATURE_THRESH_15_30": value  <= -0.00878286454826593399;
            "FEATURE_THRESH_15_31": value  <= 0.00436399597674608231;
            "FEATURE_THRESH_15_32": value  <= 0.00418047280982136726;
            "FEATURE_THRESH_15_33": value  <= -0.00045668511302210391;
            "FEATURE_THRESH_15_34": value  <= -0.00371403689496219158;
            "FEATURE_THRESH_15_35": value  <= -0.02530428953468799938;
            "FEATURE_THRESH_15_36": value  <= -0.00034454080741852522;
            "FEATURE_THRESH_15_37": value  <= -0.00083935231668874621;
            "FEATURE_THRESH_15_38": value  <= 0.01728004962205889963;
            "FEATURE_THRESH_15_39": value  <= -0.00635950779542326927;
            "FEATURE_THRESH_15_40": value  <= 0.00102981098461896181;
            "FEATURE_THRESH_15_41": value  <= 0.00101171096321195364;
            "FEATURE_THRESH_15_42": value  <= -0.01030880026519299941;
            "FEATURE_THRESH_15_43": value  <= 0.00546820182353258133;
            "FEATURE_THRESH_15_44": value  <= -0.00091696460731327534;
            "FEATURE_THRESH_15_45": value  <= 0.00239228201098740101;
            "FEATURE_THRESH_15_46": value  <= -0.00755738187581300735;
            "FEATURE_THRESH_15_47": value  <= -0.00077024032361805439;
            "FEATURE_THRESH_15_48": value  <= -0.00871259905397891998;
            "FEATURE_THRESH_15_49": value  <= -0.01030632015317680013;
            "FEATURE_THRESH_15_50": value  <= -0.00209409790113568306;
            "FEATURE_THRESH_15_51": value  <= 0.00680990517139434814;
            "FEATURE_THRESH_15_52": value  <= -0.00107460597064346075;
            "FEATURE_THRESH_15_53": value  <= 0.00215502898208796978;
            "FEATURE_THRESH_15_54": value  <= 0.03174231946468349802;
            "FEATURE_THRESH_15_55": value  <= -0.07838272303342820602;
            "FEATURE_THRESH_15_56": value  <= 0.00574151193723082542;
            "FEATURE_THRESH_15_57": value  <= -0.00290146004408597946;
            "FEATURE_THRESH_15_58": value  <= -0.00264279311522841454;
            "FEATURE_THRESH_15_59": value  <= -0.10949660092592239380;
            "FEATURE_THRESH_15_60": value  <= 0.00007407591328956187;
            "FEATURE_THRESH_15_61": value  <= -0.00050593802006915212;
            "FEATURE_THRESH_15_62": value  <= -0.00082131777890026569;
            "FEATURE_THRESH_15_63": value  <= -0.00006027653944329359;
            "FEATURE_THRESH_15_64": value  <= 0.00680651422590017319;
            "FEATURE_THRESH_15_65": value  <= 0.00172027898952364922;
            "FEATURE_THRESH_15_66": value  <= -0.00013016929733566940;
            "FEATURE_THRESH_15_67": value  <= -0.00480163889005780220;
            "FEATURE_THRESH_15_68": value  <= -0.00253993109799921513;
            "FEATURE_THRESH_15_69": value  <= -0.00142789294477552176;
            "FEATURE_THRESH_15_70": value  <= -0.02514255046844479993;
            "FEATURE_THRESH_15_71": value  <= -0.00388996093533933163;
            "FEATURE_THRESH_15_72": value  <= 0.00439474591985344887;
            "FEATURE_THRESH_15_73": value  <= 0.02467842027544980138;
            "FEATURE_THRESH_15_74": value  <= 0.03804767876863480308;
            "FEATURE_THRESH_15_75": value  <= 0.00794248655438423157;
            "FEATURE_THRESH_15_76": value  <= -0.00151100498624145985;
            "FEATURE_THRESH_15_77": value  <= 0.00642017414793372154;
            "FEATURE_THRESH_15_78": value  <= -0.00298021594062447548;
            "FEATURE_THRESH_15_79": value  <= -0.00074580078944563866;
            "FEATURE_THRESH_15_80": value  <= -0.01047095004469160082;
            "FEATURE_THRESH_15_81": value  <= 0.00933692045509815216;
            "FEATURE_THRESH_15_82": value  <= 0.02793690003454690068;
            "FEATURE_THRESH_15_83": value  <= 0.00742776785045862198;
            "FEATURE_THRESH_15_84": value  <= -0.02358450926840309839;
            "FEATURE_THRESH_15_85": value  <= 0.00114526401739567518;
            "FEATURE_THRESH_15_86": value  <= -0.00043468660442158580;
            "FEATURE_THRESH_15_87": value  <= 0.01064854022115470020;
            "FEATURE_THRESH_15_88": value  <= -0.00039418050437234342;
            "FEATURE_THRESH_15_89": value  <= -0.00013270479394122958;
            "FEATURE_THRESH_15_90": value  <= -0.00201255106367170811;
            "FEATURE_THRESH_15_91": value  <= 0.00248543196357786655;
            "FEATURE_THRESH_15_92": value  <= 0.00182378804311156273;
            "FEATURE_THRESH_15_93": value  <= -0.01665665954351430028;
            "FEATURE_THRESH_15_94": value  <= 0.00080349558265879750;
            "FEATURE_THRESH_15_95": value  <= 0.00341703789308667183;
            "FEATURE_THRESH_15_96": value  <= -0.00036222729249857366;
            "FEATURE_THRESH_15_97": value  <= -0.11630020290613170275;
            "FEATURE_THRESH_15_98": value  <= -0.01469501014798879970;
            "FEATURE_THRESH_15_99": value  <= 0.00219721300527453423;
            "FEATURE_THRESH_15_100": value  <= -0.00046965209185145795;
            "FEATURE_THRESH_15_101": value  <= 0.00651449989527463913;
            "FEATURE_THRESH_15_102": value  <= 0.02130006067454810054;
            "FEATURE_THRESH_15_103": value  <= 0.00318814092315733433;
            "FEATURE_THRESH_15_104": value  <= 0.00090019777417182922;
            "FEATURE_THRESH_15_105": value  <= -0.00517722778022289276;
            "FEATURE_THRESH_15_106": value  <= -0.00437646498903632164;
            "FEATURE_THRESH_15_107": value  <= 0.00262999604456126690;
            "FEATURE_THRESH_15_108": value  <= -0.00204586889594793320;
            "FEATURE_THRESH_15_109": value  <= 0.06948270648717880249;
            "FEATURE_THRESH_15_110": value  <= 0.02404893934726719945;
            "FEATURE_THRESH_15_111": value  <= 0.00310953403823077679;
            "FEATURE_THRESH_15_112": value  <= -0.00125032605137676001;
            "FEATURE_THRESH_15_113": value  <= -0.00102811900433152914;
            "FEATURE_THRESH_15_114": value  <= -0.00888936221599578857;
            "FEATURE_THRESH_15_115": value  <= -0.00061094801640138030;
            "FEATURE_THRESH_15_116": value  <= -0.00576863577589392662;
            "FEATURE_THRESH_15_117": value  <= 0.00185064901597797871;
            "FEATURE_THRESH_15_118": value  <= -0.09979946911334990067;
            "FEATURE_THRESH_15_119": value  <= -0.35128349065780639648;
            "FEATURE_THRESH_15_120": value  <= -0.04524457082152370108;
            "FEATURE_THRESH_15_121": value  <= 0.07148157805204390092;
            "FEATURE_THRESH_15_122": value  <= 0.00218957802280783653;
            "FEATURE_THRESH_15_123": value  <= -0.00059242651332169771;
            "FEATURE_THRESH_15_124": value  <= 0.00167883897665888071;
            "FEATURE_THRESH_15_125": value  <= -0.00221634889021515846;
            "FEATURE_THRESH_15_126": value  <= 0.00011568699846975505;
            "FEATURE_THRESH_15_127": value  <= -0.00720172887668013573;
            "FEATURE_THRESH_15_128": value  <= 0.00089081272017210722;
            "FEATURE_THRESH_15_129": value  <= 0.00019605009583756328;
            "FEATURE_THRESH_15_130": value  <= 0.00052022142335772514;
            "FEATURE_THRESH_15_131": value  <= 0.00094588572392240167;
            "FEATURE_THRESH_15_132": value  <= 0.00009169847180601211;
            "FEATURE_THRESH_15_133": value  <= 0.00218332000076770782;
            "FEATURE_THRESH_15_134": value  <= -0.00086039671441540122;
            "FEATURE_THRESH_15_135": value  <= -0.01323623955249790020;
            "FEATURE_THRESH_15_136": value  <= 0.00043376701069064438;
            "FEATURE_THRESH_16_0": value  <= -0.02484714984893799869;
            "FEATURE_THRESH_16_1": value  <= 0.00613486114889383316;
            "FEATURE_THRESH_16_2": value  <= 0.00644984981045126915;
            "FEATURE_THRESH_16_3": value  <= 0.00063491211039945483;
            "FEATURE_THRESH_16_4": value  <= 0.00140238902531564236;
            "FEATURE_THRESH_16_5": value  <= 0.00030044000595808029;
            "FEATURE_THRESH_16_6": value  <= 0.00010042409849120304;
            "FEATURE_THRESH_16_7": value  <= -0.00508414907380938530;
            "FEATURE_THRESH_16_8": value  <= -0.01953726075589659952;
            "FEATURE_THRESH_16_9": value  <= -0.00000745327406548313;
            "FEATURE_THRESH_16_10": value  <= -0.00360794598236680031;
            "FEATURE_THRESH_16_11": value  <= 0.00206975010223686695;
            "FEATURE_THRESH_16_12": value  <= -0.00046463840408250690;
            "FEATURE_THRESH_16_13": value  <= 0.00075490452582016587;
            "FEATURE_THRESH_16_14": value  <= -0.00098322238773107529;
            "FEATURE_THRESH_16_15": value  <= -0.01994064077734949980;
            "FEATURE_THRESH_16_16": value  <= 0.00376803008839488029;
            "FEATURE_THRESH_16_17": value  <= -0.00945285055786371231;
            "FEATURE_THRESH_16_18": value  <= 0.00295608490705490112;
            "FEATURE_THRESH_16_19": value  <= 0.00910787377506494522;
            "FEATURE_THRESH_16_20": value  <= 0.00182192295324057341;
            "FEATURE_THRESH_16_21": value  <= 0.01468873955309389981;
            "FEATURE_THRESH_16_22": value  <= -0.01438799034804109922;
            "FEATURE_THRESH_16_23": value  <= -0.01898664981126790136;
            "FEATURE_THRESH_16_24": value  <= 0.00115276395808905363;
            "FEATURE_THRESH_16_25": value  <= 0.01093367021530869919;
            "FEATURE_THRESH_16_26": value  <= -0.01493273023515940059;
            "FEATURE_THRESH_16_27": value  <= -0.00029970539617352188;
            "FEATURE_THRESH_16_28": value  <= 0.00416776211932301521;
            "FEATURE_THRESH_16_29": value  <= -0.00639053201302886009;
            "FEATURE_THRESH_16_30": value  <= 0.00450296094641089439;
            "FEATURE_THRESH_16_31": value  <= -0.00920403655618429184;
            "FEATURE_THRESH_16_32": value  <= 0.08132725954055790296;
            "FEATURE_THRESH_16_33": value  <= -0.15079280734062200375;
            "FEATURE_THRESH_16_34": value  <= 0.00331790093332529068;
            "FEATURE_THRESH_16_35": value  <= 0.00077402801252901554;
            "FEATURE_THRESH_16_36": value  <= 0.00068199541419744492;
            "FEATURE_THRESH_16_37": value  <= 0.00536715704947710037;
            "FEATURE_THRESH_16_38": value  <= 0.00009701866656541826;
            "FEATURE_THRESH_16_39": value  <= -0.12534089386463170834;
            "FEATURE_THRESH_16_40": value  <= -0.00525162694975733757;
            "FEATURE_THRESH_16_41": value  <= -0.00783421099185943604;
            "FEATURE_THRESH_16_42": value  <= -0.00113100698217749596;
            "FEATURE_THRESH_16_43": value  <= 0.00176011200528591871;
            "FEATURE_THRESH_16_44": value  <= -0.00081581249833106995;
            "FEATURE_THRESH_16_45": value  <= -0.00386875891126692295;
            "FEATURE_THRESH_16_46": value  <= 0.00152071297634392977;
            "FEATURE_THRESH_16_47": value  <= 0.54586738348007202148;
            "FEATURE_THRESH_16_48": value  <= 0.01565019041299819946;
            "FEATURE_THRESH_16_49": value  <= -0.01173186022788290025;
            "FEATURE_THRESH_16_50": value  <= -0.00617651222273707390;
            "FEATURE_THRESH_16_51": value  <= 0.00224576611071825027;
            "FEATURE_THRESH_16_52": value  <= -0.00519158691167831421;
            "FEATURE_THRESH_16_53": value  <= -0.02382788062095640008;
            "FEATURE_THRESH_16_54": value  <= 0.00102845800574868917;
            "FEATURE_THRESH_16_55": value  <= -0.01007885020226239985;
            "FEATURE_THRESH_16_56": value  <= 0.00261689303442835808;
            "FEATURE_THRESH_16_57": value  <= 0.00054385367548093200;
            "FEATURE_THRESH_16_58": value  <= 0.00535105122253298759;
            "FEATURE_THRESH_16_59": value  <= -0.00152747903484851122;
            "FEATURE_THRESH_16_60": value  <= -0.08062441647052759341;
            "FEATURE_THRESH_16_61": value  <= 0.02219202928245070025;
            "FEATURE_THRESH_16_62": value  <= 0.00731006311252713203;
            "FEATURE_THRESH_16_63": value  <= -0.00640630722045898438;
            "FEATURE_THRESH_16_64": value  <= -0.00076415040530264378;
            "FEATURE_THRESH_16_65": value  <= 0.00076734489994123578;
            "FEATURE_THRESH_16_66": value  <= 0.00061474501853808761;
            "FEATURE_THRESH_16_67": value  <= -0.00501052709296345711;
            "FEATURE_THRESH_16_68": value  <= -0.00869091320782899857;
            "FEATURE_THRESH_16_69": value  <= -0.01639145985245700141;
            "FEATURE_THRESH_16_70": value  <= 0.00040973909199237823;
            "FEATURE_THRESH_16_71": value  <= -0.00252422899939119816;
            "FEATURE_THRESH_16_72": value  <= 0.00050945312250405550;
            "FEATURE_THRESH_16_73": value  <= 0.00196564197540283203;
            "FEATURE_THRESH_16_74": value  <= 0.00056298897834494710;
            "FEATURE_THRESH_16_75": value  <= -0.00067946797935292125;
            "FEATURE_THRESH_16_76": value  <= 0.00728563498705625534;
            "FEATURE_THRESH_16_77": value  <= -0.01745948940515519923;
            "FEATURE_THRESH_16_78": value  <= -0.02542174980044360072;
            "FEATURE_THRESH_16_79": value  <= -0.00156476395204663277;
            "FEATURE_THRESH_16_80": value  <= 0.01144436001777649967;
            "FEATURE_THRESH_16_81": value  <= -0.00067352550104260445;
            "FEATURE_THRESH_16_82": value  <= 0.00931942090392112732;
            "FEATURE_THRESH_16_83": value  <= 0.00013328490604180843;
            "FEATURE_THRESH_16_84": value  <= -0.00788157992064952850;
            "FEATURE_THRESH_16_85": value  <= -0.00579856801778078079;
            "FEATURE_THRESH_16_86": value  <= -0.00038922499516047537;
            "FEATURE_THRESH_16_87": value  <= -0.00192886102013289928;
            "FEATURE_THRESH_16_88": value  <= 0.00842141546308994293;
            "FEATURE_THRESH_16_89": value  <= 0.00816558767110109329;
            "FEATURE_THRESH_16_90": value  <= 0.00048280550981871784;
            "FEATURE_THRESH_16_91": value  <= -0.00271866307593882084;
            "FEATURE_THRESH_16_92": value  <= -0.01250723004341129999;
            "FEATURE_THRESH_16_93": value  <= -0.02428651973605160108;
            "FEATURE_THRESH_16_94": value  <= -0.00296763307414948940;
            "FEATURE_THRESH_16_95": value  <= -0.01252899970859290037;
            "FEATURE_THRESH_16_96": value  <= -0.00101040001027286053;
            "FEATURE_THRESH_16_97": value  <= -0.00213485304266214371;
            "FEATURE_THRESH_16_98": value  <= 0.01956425979733469878;
            "FEATURE_THRESH_16_99": value  <= -0.09714634716510769930;
            "FEATURE_THRESH_16_100": value  <= 0.00450145686045289040;
            "FEATURE_THRESH_16_101": value  <= 0.00637069717049598694;
            "FEATURE_THRESH_16_102": value  <= -0.00907215289771556854;
            "FEATURE_THRESH_16_103": value  <= -0.00535372085869312286;
            "FEATURE_THRESH_16_104": value  <= -0.01093284040689469945;
            "FEATURE_THRESH_16_105": value  <= 0.00823560729622840881;
            "FEATURE_THRESH_16_106": value  <= -0.00100381602533161640;
            "FEATURE_THRESH_16_107": value  <= 0.00408591283485293388;
            "FEATURE_THRESH_16_108": value  <= 0.15485419332981109619;
            "FEATURE_THRESH_16_109": value  <= 0.00020897459762636572;
            "FEATURE_THRESH_16_110": value  <= 0.00033316991175524890;
            "FEATURE_THRESH_16_111": value  <= -0.01081340014934539968;
            "FEATURE_THRESH_16_112": value  <= 0.04565601050853729942;
            "FEATURE_THRESH_16_113": value  <= 0.00125695497263222933;
            "FEATURE_THRESH_16_114": value  <= -0.12015070021152500501;
            "FEATURE_THRESH_16_115": value  <= -0.00010533799650147557;
            "FEATURE_THRESH_16_116": value  <= -0.20703190565109250154;
            "FEATURE_THRESH_16_117": value  <= 0.00012909180077258497;
            "FEATURE_THRESH_16_118": value  <= 0.00038818528992123902;
            "FEATURE_THRESH_16_119": value  <= -0.00292436103336513042;
            "FEATURE_THRESH_16_120": value  <= 0.00083882332546636462;
            "FEATURE_THRESH_16_121": value  <= -0.00190615502651780844;
            "FEATURE_THRESH_16_122": value  <= 0.00895143486559391022;
            "FEATURE_THRESH_16_123": value  <= 0.01308345980942249992;
            "FEATURE_THRESH_16_124": value  <= -0.21159330010414120760;
            "FEATURE_THRESH_16_125": value  <= 0.00314932502806186676;
            "FEATURE_THRESH_16_126": value  <= 0.00039754100725986063;
            "FEATURE_THRESH_16_127": value  <= -0.00138144800439476967;
            "FEATURE_THRESH_16_128": value  <= -0.00058122188784182072;
            "FEATURE_THRESH_16_129": value  <= -0.00239053298719227314;
            "FEATURE_THRESH_16_130": value  <= 0.02726892940700050005;
            "FEATURE_THRESH_16_131": value  <= -0.00376583589240908623;
            "FEATURE_THRESH_16_132": value  <= -0.00149034895002841949;
            "FEATURE_THRESH_16_133": value  <= -0.01742823049426079837;
            "FEATURE_THRESH_16_134": value  <= -0.01527803018689159915;
            "FEATURE_THRESH_16_135": value  <= 0.03199560940265659681;
            "FEATURE_THRESH_16_136": value  <= -0.00382567103952169418;
            "FEATURE_THRESH_16_137": value  <= -0.00851864367723464966;
            "FEATURE_THRESH_16_138": value  <= 0.00090641621500253677;
            "FEATURE_THRESH_16_139": value  <= 0.01034484989941119974;
            "FEATURE_THRESH_17_0": value  <= 0.00789818260818719864;
            "FEATURE_THRESH_17_1": value  <= 0.00161701603792607784;
            "FEATURE_THRESH_17_2": value  <= -0.00055449741194024682;
            "FEATURE_THRESH_17_3": value  <= 0.00154289801139384508;
            "FEATURE_THRESH_17_4": value  <= -0.00103294500149786472;
            "FEATURE_THRESH_17_5": value  <= 0.00077698158565908670;
            "FEATURE_THRESH_17_6": value  <= 0.14320300519466400146;
            "FEATURE_THRESH_17_7": value  <= -0.00738664902746677399;
            "FEATURE_THRESH_17_8": value  <= -0.00062936742324382067;
            "FEATURE_THRESH_17_9": value  <= 0.00078893528552725911;
            "FEATURE_THRESH_17_10": value  <= -0.01222805026918650020;
            "FEATURE_THRESH_17_11": value  <= 0.00354202394373714924;
            "FEATURE_THRESH_17_12": value  <= -0.00105853204149752855;
            "FEATURE_THRESH_17_13": value  <= 0.00001493566014687531;
            "FEATURE_THRESH_17_14": value  <= 0.00525377085432410240;
            "FEATURE_THRESH_17_15": value  <= -0.00823380239307880402;
            "FEATURE_THRESH_17_16": value  <= 0.00002186681012972258;
            "FEATURE_THRESH_17_17": value  <= -0.00381502299569547176;
            "FEATURE_THRESH_17_18": value  <= 0.00111058796755969524;
            "FEATURE_THRESH_17_19": value  <= -0.00577076897025108337;
            "FEATURE_THRESH_17_20": value  <= -0.00301583390682935715;
            "FEATURE_THRESH_17_21": value  <= -0.00085453689098358154;
            "FEATURE_THRESH_17_22": value  <= 0.01105051022022959968;
            "FEATURE_THRESH_17_23": value  <= 0.04260583966970440256;
            "FEATURE_THRESH_17_24": value  <= -0.00307817501015961170;
            "FEATURE_THRESH_17_25": value  <= -0.00548157282173633575;
            "FEATURE_THRESH_17_26": value  <= 0.00318818609230220318;
            "FEATURE_THRESH_17_27": value  <= 0.00035947180003859103;
            "FEATURE_THRESH_17_28": value  <= -0.00407050317153334618;
            "FEATURE_THRESH_17_29": value  <= -0.01459417026489969946;
            "FEATURE_THRESH_17_30": value  <= -0.00011947689927183092;
            "FEATURE_THRESH_17_31": value  <= -0.00069344649091362953;
            "FEATURE_THRESH_17_32": value  <= 0.00001483479991293280;
            "FEATURE_THRESH_17_33": value  <= 0.00902969855815172195;
            "FEATURE_THRESH_17_34": value  <= -0.00806408189237117767;
            "FEATURE_THRESH_17_35": value  <= 0.02606211975216870050;
            "FEATURE_THRESH_17_36": value  <= 0.01731465943157670107;
            "FEATURE_THRESH_17_37": value  <= 0.02266664057970050120;
            "FEATURE_THRESH_17_38": value  <= -0.00219659297727048397;
            "FEATURE_THRESH_17_39": value  <= -0.00952824763953685760;
            "FEATURE_THRESH_17_40": value  <= 0.00809436198323965073;
            "FEATURE_THRESH_17_41": value  <= -0.07287733256816859850;
            "FEATURE_THRESH_17_42": value  <= -0.00690095219761133194;
            "FEATURE_THRESH_17_43": value  <= -0.01130823977291580025;
            "FEATURE_THRESH_17_44": value  <= 0.05961320176720619896;
            "FEATURE_THRESH_17_45": value  <= -0.00286246207542717457;
            "FEATURE_THRESH_17_46": value  <= 0.00447814492508769035;
            "FEATURE_THRESH_17_47": value  <= -0.00175132404547184706;
            "FEATURE_THRESH_17_48": value  <= 0.04016342014074329725;
            "FEATURE_THRESH_17_49": value  <= 0.00034768949262797832;
            "FEATURE_THRESH_17_50": value  <= 0.00265516503714025021;
            "FEATURE_THRESH_17_51": value  <= -0.00877062790095806122;
            "FEATURE_THRESH_17_52": value  <= -0.00551220914348959923;
            "FEATURE_THRESH_17_53": value  <= 0.00068672042107209563;
            "FEATURE_THRESH_17_54": value  <= 0.00056019669864326715;
            "FEATURE_THRESH_17_55": value  <= 0.00241437694057822227;
            "FEATURE_THRESH_17_56": value  <= -0.00156809005420655012;
            "FEATURE_THRESH_17_57": value  <= -0.00368274911306798458;
            "FEATURE_THRESH_17_58": value  <= -0.00029409190756268799;
            "FEATURE_THRESH_17_59": value  <= 0.00042847759323194623;
            "FEATURE_THRESH_17_60": value  <= -0.00488170702010393143;
            "FEATURE_THRESH_17_61": value  <= 0.00027272020815871656;
            "FEATURE_THRESH_17_62": value  <= 0.00020947199664078653;
            "FEATURE_THRESH_17_63": value  <= 0.04850118979811669784;
            "FEATURE_THRESH_17_64": value  <= -0.00451664114370942116;
            "FEATURE_THRESH_17_65": value  <= -0.01229168009012939974;
            "FEATURE_THRESH_17_66": value  <= 0.00048549679922871292;
            "FEATURE_THRESH_17_67": value  <= 0.03055604919791219884;
            "FEATURE_THRESH_17_68": value  <= -0.00015105320198927075;
            "FEATURE_THRESH_17_69": value  <= 0.00249374401755630970;
            "FEATURE_THRESH_17_70": value  <= -0.01238213013857599951;
            "FEATURE_THRESH_17_71": value  <= -0.00513334618881344795;
            "FEATURE_THRESH_17_72": value  <= 0.00051919277757406235;
            "FEATURE_THRESH_17_73": value  <= 0.15060420334339139070;
            "FEATURE_THRESH_17_74": value  <= 0.00771441496908664703;
            "FEATURE_THRESH_17_75": value  <= 0.00944435223937034607;
            "FEATURE_THRESH_17_76": value  <= 0.00025006249779835343;
            "FEATURE_THRESH_17_77": value  <= -0.00330771505832672119;
            "FEATURE_THRESH_17_78": value  <= 0.00074048910755664110;
            "FEATURE_THRESH_17_79": value  <= 0.04409205168485640092;
            "FEATURE_THRESH_17_80": value  <= 0.00336399092338979244;
            "FEATURE_THRESH_17_81": value  <= -0.00397600792348384857;
            "FEATURE_THRESH_17_82": value  <= 0.00277169304899871349;
            "FEATURE_THRESH_17_83": value  <= -0.00024123019829858094;
            "FEATURE_THRESH_17_84": value  <= 0.00049425667384639382;
            "FEATURE_THRESH_17_85": value  <= -0.00038876468897797167;
            "FEATURE_THRESH_17_86": value  <= -0.05004889890551569853;
            "FEATURE_THRESH_17_87": value  <= -0.03663548082113270155;
            "FEATURE_THRESH_17_88": value  <= 0.00242735794745385647;
            "FEATURE_THRESH_17_89": value  <= 0.00195580301806330681;
            "FEATURE_THRESH_17_90": value  <= -0.00174946105107665062;
            "FEATURE_THRESH_17_91": value  <= 0.01395507995039219941;
            "FEATURE_THRESH_17_92": value  <= -0.00021896739781368524;
            "FEATURE_THRESH_17_93": value  <= -0.00151313096284866333;
            "FEATURE_THRESH_17_94": value  <= -0.00436228001490235329;
            "FEATURE_THRESH_17_95": value  <= 0.06516058743000030518;
            "FEATURE_THRESH_17_96": value  <= -0.00235673994757235050;
            "FEATURE_THRESH_17_97": value  <= 0.01514665968716140051;
            "FEATURE_THRESH_17_98": value  <= -0.02285096049308779978;
            "FEATURE_THRESH_17_99": value  <= 0.00488676503300666809;
            "FEATURE_THRESH_17_100": value  <= 0.00176195998210459948;
            "FEATURE_THRESH_17_101": value  <= -0.00129425199702382088;
            "FEATURE_THRESH_17_102": value  <= 0.01092994958162309994;
            "FEATURE_THRESH_17_103": value  <= 0.00002995848990394734;
            "FEATURE_THRESH_17_104": value  <= -0.00658843619748950005;
            "FEATURE_THRESH_17_105": value  <= 0.00325277796946465969;
            "FEATURE_THRESH_17_106": value  <= -0.00404357397928833961;
            "FEATURE_THRESH_17_107": value  <= -0.00125235400628298521;
            "FEATURE_THRESH_17_108": value  <= 0.00019246719602961093;
            "FEATURE_THRESH_17_109": value  <= -0.03858967125415799920;
            "FEATURE_THRESH_17_110": value  <= 0.00015489870565943420;
            "FEATURE_THRESH_17_111": value  <= -0.03376384824514389732;
            "FEATURE_THRESH_17_112": value  <= -0.00826570671051740646;
            "FEATURE_THRESH_17_113": value  <= 0.00001448144030291587;
            "FEATURE_THRESH_17_114": value  <= 0.00001495129981776700;
            "FEATURE_THRESH_17_115": value  <= -0.01874179951846599926;
            "FEATURE_THRESH_17_116": value  <= 0.00175722397398203611;
            "FEATURE_THRESH_17_117": value  <= -0.00313911191187798977;
            "FEATURE_THRESH_17_118": value  <= 0.00006665677938144654;
            "FEATURE_THRESH_17_119": value  <= 0.00677434215322136879;
            "FEATURE_THRESH_17_120": value  <= -0.00738681619986891747;
            "FEATURE_THRESH_17_121": value  <= 0.01404093019664289996;
            "FEATURE_THRESH_17_122": value  <= -0.00552583299577236176;
            "FEATURE_THRESH_17_123": value  <= 0.38684239983558660336;
            "FEATURE_THRESH_17_124": value  <= 0.00011459240340627730;
            "FEATURE_THRESH_17_125": value  <= -0.01846756972372530156;
            "FEATURE_THRESH_17_126": value  <= -0.00045907011372037232;
            "FEATURE_THRESH_17_127": value  <= 0.00125275400932878256;
            "FEATURE_THRESH_17_128": value  <= 0.00149106094613671303;
            "FEATURE_THRESH_17_129": value  <= -0.00075435562757775187;
            "FEATURE_THRESH_17_130": value  <= -0.00694788387045264244;
            "FEATURE_THRESH_17_131": value  <= 0.00028092920547351241;
            "FEATURE_THRESH_17_132": value  <= 0.00096073717577382922;
            "FEATURE_THRESH_17_133": value  <= -0.00026883929967880249;
            "FEATURE_THRESH_17_134": value  <= 0.00215993705205619335;
            "FEATURE_THRESH_17_135": value  <= 0.00562353013083338737;
            "FEATURE_THRESH_17_136": value  <= -0.00502439914271235466;
            "FEATURE_THRESH_17_137": value  <= -0.00976116396486759186;
            "FEATURE_THRESH_17_138": value  <= 0.00415151007473468781;
            "FEATURE_THRESH_17_139": value  <= 0.00624650809913873672;
            "FEATURE_THRESH_17_140": value  <= -0.00705974781885743141;
            "FEATURE_THRESH_17_141": value  <= -0.00205877097323536873;
            "FEATURE_THRESH_17_142": value  <= -0.00241460604593157768;
            "FEATURE_THRESH_17_143": value  <= -0.00148176099173724651;
            "FEATURE_THRESH_17_144": value  <= -0.00630164006724953651;
            "FEATURE_THRESH_17_145": value  <= 0.00347634288482367992;
            "FEATURE_THRESH_17_146": value  <= -0.02225087024271489924;
            "FEATURE_THRESH_17_147": value  <= -0.03061255067586899845;
            "FEATURE_THRESH_17_148": value  <= 0.01305747963488100051;
            "FEATURE_THRESH_17_149": value  <= -0.00060095742810517550;
            "FEATURE_THRESH_17_150": value  <= -0.00041514250915497541;
            "FEATURE_THRESH_17_151": value  <= -0.01377629023045300050;
            "FEATURE_THRESH_17_152": value  <= -0.03229650855064390008;
            "FEATURE_THRESH_17_153": value  <= 0.05355697870254520071;
            "FEATURE_THRESH_17_154": value  <= 0.00818895455449819565;
            "FEATURE_THRESH_17_155": value  <= 0.00021055320394225419;
            "FEATURE_THRESH_17_156": value  <= -0.00243827304802834988;
            "FEATURE_THRESH_17_157": value  <= 0.00328355701640248299;
            "FEATURE_THRESH_17_158": value  <= 0.00237295706756412983;
            "FEATURE_THRESH_17_159": value  <= -0.00145416997838765383;
            "FEATURE_THRESH_18_0": value  <= 0.05575523898005489698;
            "FEATURE_THRESH_18_1": value  <= 0.00247302488423883915;
            "FEATURE_THRESH_18_2": value  <= -0.00035031698644161224;
            "FEATURE_THRESH_18_3": value  <= 0.00054167630150914192;
            "FEATURE_THRESH_18_4": value  <= 0.00077193678589537740;
            "FEATURE_THRESH_18_5": value  <= -0.00159992196131497622;
            "FEATURE_THRESH_18_6": value  <= -0.00011832080053864047;
            "FEATURE_THRESH_18_7": value  <= 0.00032909031142480671;
            "FEATURE_THRESH_18_8": value  <= 0.00029518108931370080;
            "FEATURE_THRESH_18_9": value  <= 0.00009046671038959177;
            "FEATURE_THRESH_18_10": value  <= 0.00001500719008618035;
            "FEATURE_THRESH_18_11": value  <= 0.13935610651969909668;
            "FEATURE_THRESH_18_12": value  <= 0.00164619903080165386;
            "FEATURE_THRESH_18_13": value  <= 0.00049984431825578213;
            "FEATURE_THRESH_18_14": value  <= -0.00109712802805006504;
            "FEATURE_THRESH_18_15": value  <= 0.00066919892560690641;
            "FEATURE_THRESH_18_16": value  <= 0.00086471042595803738;
            "FEATURE_THRESH_18_17": value  <= -0.00027182599296793342;
            "FEATURE_THRESH_18_18": value  <= 0.00003024949910468422;
            "FEATURE_THRESH_18_19": value  <= -0.00852258969098329544;
            "FEATURE_THRESH_18_20": value  <= 0.00167055602651089430;
            "FEATURE_THRESH_18_21": value  <= -0.00714338384568691254;
            "FEATURE_THRESH_18_22": value  <= -0.01631936989724639894;
            "FEATURE_THRESH_18_23": value  <= 0.00480342609807848930;
            "FEATURE_THRESH_18_24": value  <= -0.00754219293594360352;
            "FEATURE_THRESH_18_25": value  <= -0.01436311006546019987;
            "FEATURE_THRESH_18_26": value  <= 0.00089063588529825211;
            "FEATURE_THRESH_18_27": value  <= -0.00440601911395788193;
            "FEATURE_THRESH_18_28": value  <= -0.00018862540309783071;
            "FEATURE_THRESH_18_29": value  <= -0.00379792810417711735;
            "FEATURE_THRESH_18_30": value  <= 0.00014627049677073956;
            "FEATURE_THRESH_18_31": value  <= -0.00004916463876725175;
            "FEATURE_THRESH_18_32": value  <= -0.03358250111341479910;
            "FEATURE_THRESH_18_33": value  <= -0.00353393098339438438;
            "FEATURE_THRESH_18_34": value  <= 0.00501441117376089096;
            "FEATURE_THRESH_18_35": value  <= 0.01881737075746060112;
            "FEATURE_THRESH_18_36": value  <= -0.00134343397803604603;
            "FEATURE_THRESH_18_37": value  <= 0.00175579602364450693;
            "FEATURE_THRESH_18_38": value  <= -0.09563746303319929642;
            "FEATURE_THRESH_18_39": value  <= -0.02224122919142250063;
            "FEATURE_THRESH_18_40": value  <= -0.01557581964880229951;
            "FEATURE_THRESH_18_41": value  <= 0.00535991182550787926;
            "FEATURE_THRESH_18_42": value  <= -0.02176349982619290094;
            "FEATURE_THRESH_18_43": value  <= -0.16561590135097500887;
            "FEATURE_THRESH_18_44": value  <= 0.00016461320046801120;
            "FEATURE_THRESH_18_45": value  <= -0.00890775024890899658;
            "FEATURE_THRESH_18_46": value  <= 0.00086346449097618461;
            "FEATURE_THRESH_18_47": value  <= -0.00137517601251602173;
            "FEATURE_THRESH_18_48": value  <= -0.00140812399331480265;
            "FEATURE_THRESH_18_49": value  <= -0.00393428886309266090;
            "FEATURE_THRESH_18_50": value  <= -0.03196692839264869690;
            "FEATURE_THRESH_18_51": value  <= -0.00001508928016846767;
            "FEATURE_THRESH_18_52": value  <= 0.00051994470413774252;
            "FEATURE_THRESH_18_53": value  <= -0.00342204608023166656;
            "FEATURE_THRESH_18_54": value  <= 0.00017723299970384687;
            "FEATURE_THRESH_18_55": value  <= 0.00157167599536478519;
            "FEATURE_THRESH_18_56": value  <= -0.00890413299202919006;
            "FEATURE_THRESH_18_57": value  <= 0.00040677518700249493;
            "FEATURE_THRESH_18_58": value  <= 0.00676047801971435547;
            "FEATURE_THRESH_18_59": value  <= 0.00291000888682901859;
            "FEATURE_THRESH_18_60": value  <= 0.00138854596298187971;
            "FEATURE_THRESH_18_61": value  <= -0.07676426321268080277;
            "FEATURE_THRESH_18_62": value  <= -0.00022688310127705336;
            "FEATURE_THRESH_18_63": value  <= -0.00630941521376371384;
            "FEATURE_THRESH_18_64": value  <= -0.11007279902696609497;
            "FEATURE_THRESH_18_65": value  <= 0.00028619659133255482;
            "FEATURE_THRESH_18_66": value  <= 0.00002942532955785282;
            "FEATURE_THRESH_18_67": value  <= -0.02488657087087629838;
            "FEATURE_THRESH_18_68": value  <= 0.03314885124564170144;
            "FEATURE_THRESH_18_69": value  <= 0.00078491691965609789;
            "FEATURE_THRESH_18_70": value  <= 0.00470871897414326668;
            "FEATURE_THRESH_18_71": value  <= 0.00241444795392453671;
            "FEATURE_THRESH_18_72": value  <= 0.00195231800898909569;
            "FEATURE_THRESH_18_73": value  <= 0.00130319804884493351;
            "FEATURE_THRESH_18_74": value  <= 0.00447354977950453758;
            "FEATURE_THRESH_18_75": value  <= -0.00266528688371181488;
            "FEATURE_THRESH_18_76": value  <= 0.00013666770246345550;
            "FEATURE_THRESH_18_77": value  <= -0.01712645031511780130;
            "FEATURE_THRESH_18_78": value  <= -0.00026601430727168918;
            "FEATURE_THRESH_18_79": value  <= -0.02293238043785100072;
            "FEATURE_THRESH_18_80": value  <= 0.00233165500685572624;
            "FEATURE_THRESH_18_81": value  <= 0.01692566089332099913;
            "FEATURE_THRESH_18_82": value  <= -0.00898588262498378754;
            "FEATURE_THRESH_18_83": value  <= -0.01187469996511940004;
            "FEATURE_THRESH_18_84": value  <= 0.00019350569345988333;
            "FEATURE_THRESH_18_85": value  <= 0.00587134901434183121;
            "FEATURE_THRESH_18_86": value  <= -0.24838790297508239746;
            "FEATURE_THRESH_18_87": value  <= 0.01225600019097329921;
            "FEATURE_THRESH_18_88": value  <= 0.00083990179700776935;
            "FEATURE_THRESH_18_89": value  <= 0.00254073692485690117;
            "FEATURE_THRESH_18_90": value  <= -0.01482242997735739969;
            "FEATURE_THRESH_18_91": value  <= -0.00579739594832062721;
            "FEATURE_THRESH_18_92": value  <= 0.00072662148158997297;
            "FEATURE_THRESH_18_93": value  <= -0.01723258011043070012;
            "FEATURE_THRESH_18_94": value  <= 0.00786240864545106888;
            "FEATURE_THRESH_18_95": value  <= -0.00473436200991272926;
            "FEATURE_THRESH_18_96": value  <= 0.00083048478700220585;
            "FEATURE_THRESH_18_97": value  <= 0.00766021991148591042;
            "FEATURE_THRESH_18_98": value  <= -0.00410483777523040771;
            "FEATURE_THRESH_18_99": value  <= 0.00485125789418816566;
            "FEATURE_THRESH_18_100": value  <= 0.00099896453320980072;
            "FEATURE_THRESH_18_101": value  <= -0.27023631334304809570;
            "FEATURE_THRESH_18_102": value  <= -0.01309068035334350066;
            "FEATURE_THRESH_18_103": value  <= -0.00943427905440330505;
            "FEATURE_THRESH_18_104": value  <= -0.00154820398893207312;
            "FEATURE_THRESH_18_105": value  <= 0.00537461321800947189;
            "FEATURE_THRESH_18_106": value  <= 0.00157867697998881340;
            "FEATURE_THRESH_18_107": value  <= 0.00368560501374304295;
            "FEATURE_THRESH_18_108": value  <= 0.00938870199024677277;
            "FEATURE_THRESH_18_109": value  <= 0.01279263012111189930;
            "FEATURE_THRESH_18_110": value  <= -0.00336610409431159496;
            "FEATURE_THRESH_18_111": value  <= 0.00039771420415490866;
            "FEATURE_THRESH_18_112": value  <= 0.00148680305574089289;
            "FEATURE_THRESH_18_113": value  <= -0.08868674933910369873;
            "FEATURE_THRESH_18_114": value  <= -0.00007429611287079751;
            "FEATURE_THRESH_18_115": value  <= -0.00001493293984822231;
            "FEATURE_THRESH_18_116": value  <= 0.00591622386127710342;
            "FEATURE_THRESH_18_117": value  <= 0.00111416401341557503;
            "FEATURE_THRESH_18_118": value  <= 0.00008924936264520512;
            "FEATURE_THRESH_18_119": value  <= 0.00253195106051862240;
            "FEATURE_THRESH_18_120": value  <= 0.01242620032280680048;
            "FEATURE_THRESH_18_121": value  <= 0.02833575010299679842;
            "FEATURE_THRESH_18_122": value  <= 0.00661658821627497673;
            "FEATURE_THRESH_18_123": value  <= 0.00804687663912773132;
            "FEATURE_THRESH_18_124": value  <= -0.00111939804628491402;
            "FEATURE_THRESH_18_125": value  <= 0.01327759027481079969;
            "FEATURE_THRESH_18_126": value  <= 0.00048794739996083081;
            "FEATURE_THRESH_18_127": value  <= 0.01124317012727260069;
            "FEATURE_THRESH_18_128": value  <= -0.00089896668214350939;
            "FEATURE_THRESH_18_129": value  <= 0.00666771596297621727;
            "FEATURE_THRESH_18_130": value  <= 0.02894729934632779902;
            "FEATURE_THRESH_18_131": value  <= -0.02340004965662960054;
            "FEATURE_THRESH_18_132": value  <= -0.08911705017089839587;
            "FEATURE_THRESH_18_133": value  <= -0.01405460014939310075;
            "FEATURE_THRESH_18_134": value  <= 0.00812393985688686371;
            "FEATURE_THRESH_18_135": value  <= -0.00499646505340933800;
            "FEATURE_THRESH_18_136": value  <= 0.00312539702281355858;
            "FEATURE_THRESH_18_137": value  <= 0.00676696421578526497;
            "FEATURE_THRESH_18_138": value  <= -0.00237114401534199715;
            "FEATURE_THRESH_18_139": value  <= -0.00535227917134761810;
            "FEATURE_THRESH_18_140": value  <= -0.01596885919570920076;
            "FEATURE_THRESH_18_141": value  <= 0.00476760603487491608;
            "FEATURE_THRESH_18_142": value  <= -0.00247146910987794399;
            "FEATURE_THRESH_18_143": value  <= -0.00071033788844943047;
            "FEATURE_THRESH_18_144": value  <= -0.14117559790611269865;
            "FEATURE_THRESH_18_145": value  <= 0.10651809722185140439;
            "FEATURE_THRESH_18_146": value  <= -0.05274474993348120255;
            "FEATURE_THRESH_18_147": value  <= -0.00474317604675889015;
            "FEATURE_THRESH_18_148": value  <= 0.00099676765967160463;
            "FEATURE_THRESH_18_149": value  <= 0.00802841316908597946;
            "FEATURE_THRESH_18_150": value  <= 0.00086025858763605356;
            "FEATURE_THRESH_18_151": value  <= 0.00093191501218825579;
            "FEATURE_THRESH_18_152": value  <= -0.00250820606015622616;
            "FEATURE_THRESH_18_153": value  <= -0.00213787611573934555;
            "FEATURE_THRESH_18_154": value  <= -0.00215460499748587608;
            "FEATURE_THRESH_18_155": value  <= -0.00762140098959207535;
            "FEATURE_THRESH_18_156": value  <= 0.00220553600229322910;
            "FEATURE_THRESH_18_157": value  <= 0.00125869503244757652;
            "FEATURE_THRESH_18_158": value  <= -0.00509267207235097885;
            "FEATURE_THRESH_18_159": value  <= -0.00250957394018769264;
            "FEATURE_THRESH_18_160": value  <= -0.07732755690813060412;
            "FEATURE_THRESH_18_161": value  <= -0.04148581996560100210;
            "FEATURE_THRESH_18_162": value  <= 0.00010355669655837119;
            "FEATURE_THRESH_18_163": value  <= 0.00132558098994195461;
            "FEATURE_THRESH_18_164": value  <= -0.00805987324565649033;
            "FEATURE_THRESH_18_165": value  <= 0.01905862055718900161;
            "FEATURE_THRESH_18_166": value  <= -0.03505789116024970314;
            "FEATURE_THRESH_18_167": value  <= 0.00572960590943694115;
            "FEATURE_THRESH_18_168": value  <= -0.01164832990616559982;
            "FEATURE_THRESH_18_169": value  <= 0.00145444797817617655;
            "FEATURE_THRESH_18_170": value  <= -0.00025030909455381334;
            "FEATURE_THRESH_18_171": value  <= -0.00082907272735610604;
            "FEATURE_THRESH_18_172": value  <= 0.00108622096013277769;
            "FEATURE_THRESH_18_173": value  <= 0.00020000500080641359;
            "FEATURE_THRESH_18_174": value  <= 0.00292129209265112877;
            "FEATURE_THRESH_18_175": value  <= 0.02538740076124669856;
            "FEATURE_THRESH_18_176": value  <= -0.00319684692658483982;
            "FEATURE_THRESH_19_0": value  <= 0.00580317387357354164;
            "FEATURE_THRESH_19_1": value  <= -0.00900030694901943207;
            "FEATURE_THRESH_19_2": value  <= -0.00115496595390141010;
            "FEATURE_THRESH_19_3": value  <= -0.00110698502976447344;
            "FEATURE_THRESH_19_4": value  <= 0.00010308309720130637;
            "FEATURE_THRESH_19_5": value  <= -0.00509848399087786674;
            "FEATURE_THRESH_19_6": value  <= 0.00082572200335562229;
            "FEATURE_THRESH_19_7": value  <= 0.00997833255678415298;
            "FEATURE_THRESH_19_8": value  <= -0.03740252926945689810;
            "FEATURE_THRESH_19_9": value  <= 0.00485482579097151756;
            "FEATURE_THRESH_19_10": value  <= -0.00186644704081118107;
            "FEATURE_THRESH_19_11": value  <= 0.01688889041543010019;
            "FEATURE_THRESH_19_12": value  <= -0.00583726214244961739;
            "FEATURE_THRESH_19_13": value  <= -0.00147137395106256008;
            "FEATURE_THRESH_19_14": value  <= -0.00115229503717273474;
            "FEATURE_THRESH_19_15": value  <= -0.00425603007897734642;
            "FEATURE_THRESH_19_16": value  <= -0.00673782918602228165;
            "FEATURE_THRESH_19_17": value  <= 0.01138267014175649988;
            "FEATURE_THRESH_19_18": value  <= 0.00517947087064385414;
            "FEATURE_THRESH_19_19": value  <= -0.11743789911270140214;
            "FEATURE_THRESH_19_20": value  <= 0.02870344929397109987;
            "FEATURE_THRESH_19_21": value  <= 0.00482310308143496513;
            "FEATURE_THRESH_19_22": value  <= 0.00267985300160944462;
            "FEATURE_THRESH_19_23": value  <= 0.00805040821433067322;
            "FEATURE_THRESH_19_24": value  <= 0.00480549596250057220;
            "FEATURE_THRESH_19_25": value  <= -0.00224201590754091740;
            "FEATURE_THRESH_19_26": value  <= -0.01375771034508939915;
            "FEATURE_THRESH_19_27": value  <= -0.10338299721479420057;
            "FEATURE_THRESH_19_28": value  <= -0.00944320857524871826;
            "FEATURE_THRESH_19_29": value  <= 0.00080271181650459766;
            "FEATURE_THRESH_19_30": value  <= -0.00419456698000431061;
            "FEATURE_THRESH_19_31": value  <= 0.01094221044331790058;
            "FEATURE_THRESH_19_32": value  <= -0.00057841069065034389;
            "FEATURE_THRESH_19_33": value  <= -0.00208886200562119484;
            "FEATURE_THRESH_19_34": value  <= 0.00323839695192873478;
            "FEATURE_THRESH_19_35": value  <= 0.00490750279277563095;
            "FEATURE_THRESH_19_36": value  <= -0.03227794170379640060;
            "FEATURE_THRESH_19_37": value  <= -0.00897112302482128143;
            "FEATURE_THRESH_19_38": value  <= 0.01532108988612890070;
            "FEATURE_THRESH_19_39": value  <= 0.00208555697463452816;
            "FEATURE_THRESH_19_40": value  <= 0.00506150210276246071;
            "FEATURE_THRESH_19_41": value  <= -0.00371747510507702827;
            "FEATURE_THRESH_19_42": value  <= -0.01217050012201069918;
            "FEATURE_THRESH_19_43": value  <= 0.00462483987212181091;
            "FEATURE_THRESH_19_44": value  <= -0.00021040429419372231;
            "FEATURE_THRESH_19_45": value  <= -0.01464178040623659999;
            "FEATURE_THRESH_19_46": value  <= 0.00331994891166687012;
            "FEATURE_THRESH_19_47": value  <= 0.00372368795797228813;
            "FEATURE_THRESH_19_48": value  <= 0.00082951161311939359;
            "FEATURE_THRESH_19_49": value  <= -0.01140849012881520012;
            "FEATURE_THRESH_19_50": value  <= -0.00453201215714216232;
            "FEATURE_THRESH_19_51": value  <= 0.00512760179117321968;
            "FEATURE_THRESH_19_52": value  <= 0.00985831581056118011;
            "FEATURE_THRESH_19_53": value  <= 0.03698591887950899992;
            "FEATURE_THRESH_19_54": value  <= 0.00464911619201302528;
            "FEATURE_THRESH_19_55": value  <= -0.00426647020503878593;
            "FEATURE_THRESH_19_56": value  <= -0.00047956590424291790;
            "FEATURE_THRESH_19_57": value  <= 0.00368271605111658573;
            "FEATURE_THRESH_19_58": value  <= -0.01005988009274010053;
            "FEATURE_THRESH_19_59": value  <= -0.00030361840617842972;
            "FEATURE_THRESH_19_60": value  <= -0.00145454797893762589;
            "FEATURE_THRESH_19_61": value  <= 0.00165152095723897219;
            "FEATURE_THRESH_19_62": value  <= -0.00784686394035816193;
            "FEATURE_THRESH_19_63": value  <= -0.00512598501518368721;
            "FEATURE_THRESH_19_64": value  <= -0.03689096122980119880;
            "FEATURE_THRESH_19_65": value  <= 0.00024035639944486320;
            "FEATURE_THRESH_19_66": value  <= -0.00001515016992925666;
            "FEATURE_THRESH_19_67": value  <= 0.00221084710210561752;
            "FEATURE_THRESH_19_68": value  <= -0.00115686201024800539;
            "FEATURE_THRESH_19_69": value  <= 0.00499962922185659409;
            "FEATURE_THRESH_19_70": value  <= -0.00146561895962804556;
            "FEATURE_THRESH_19_71": value  <= -0.00119750399608165026;
            "FEATURE_THRESH_19_72": value  <= -0.00449543306604027748;
            "FEATURE_THRESH_19_73": value  <= 0.00014997160178609192;
            "FEATURE_THRESH_19_74": value  <= 0.00263915094546973705;
            "FEATURE_THRESH_19_75": value  <= -0.00029368131072260439;
            "FEATURE_THRESH_19_76": value  <= 0.00142117601353675127;
            "FEATURE_THRESH_19_77": value  <= 0.07942763715982439909;
            "FEATURE_THRESH_19_78": value  <= 0.07993750274181370130;
            "FEATURE_THRESH_19_79": value  <= 0.01108925975859170049;
            "FEATURE_THRESH_19_80": value  <= 0.00016560709627810866;
            "FEATURE_THRESH_19_81": value  <= -0.00533542921766638756;
            "FEATURE_THRESH_19_82": value  <= 0.00112872605677694082;
            "FEATURE_THRESH_19_83": value  <= -0.02196921966969970011;
            "FEATURE_THRESH_19_84": value  <= -0.00021775320055894554;
            "FEATURE_THRESH_19_85": value  <= 0.00020200149447191507;
            "FEATURE_THRESH_19_86": value  <= -0.02173314988613130050;
            "FEATURE_THRESH_19_87": value  <= -0.00084399932529777288;
            "FEATURE_THRESH_19_88": value  <= -0.00043895249837078154;
            "FEATURE_THRESH_19_89": value  <= 0.00150924001354724169;
            "FEATURE_THRESH_19_90": value  <= -0.00355478399433195591;
            "FEATURE_THRESH_19_91": value  <= 0.00048191400128416717;
            "FEATURE_THRESH_19_92": value  <= -0.00602643983438611031;
            "FEATURE_THRESH_19_93": value  <= -0.01166814006865020056;
            "FEATURE_THRESH_19_94": value  <= -0.00287183700129389763;
            "FEATURE_THRESH_19_95": value  <= 0.01705116964876650029;
            "FEATURE_THRESH_19_96": value  <= -0.01335208024829630073;
            "FEATURE_THRESH_19_97": value  <= -0.00039301801007241011;
            "FEATURE_THRESH_19_98": value  <= 0.00304833496920764446;
            "FEATURE_THRESH_19_99": value  <= -0.00435792887583374977;
            "FEATURE_THRESH_19_100": value  <= 0.00566610181704163551;
            "FEATURE_THRESH_19_101": value  <= 0.00006067733920644969;
            "FEATURE_THRESH_19_102": value  <= 0.03673816099762920034;
            "FEATURE_THRESH_19_103": value  <= 0.00865281373262405396;
            "FEATURE_THRESH_19_104": value  <= -0.15371359884738919344;
            "FEATURE_THRESH_19_105": value  <= -0.00041560421232134104;
            "FEATURE_THRESH_19_106": value  <= -0.00126401695888489485;
            "FEATURE_THRESH_19_107": value  <= -0.00354733411222696304;
            "FEATURE_THRESH_19_108": value  <= 0.00003001906952704303;
            "FEATURE_THRESH_19_109": value  <= 0.00131130195222795010;
            "FEATURE_THRESH_19_110": value  <= -0.00133747095242142677;
            "FEATURE_THRESH_19_111": value  <= 0.02087670937180520145;
            "FEATURE_THRESH_19_112": value  <= -0.00754979485645890236;
            "FEATURE_THRESH_19_113": value  <= 0.02418855018913750043;
            "FEATURE_THRESH_19_114": value  <= -0.00293588289059698582;
            "FEATURE_THRESH_19_115": value  <= 0.05755792930722240103;
            "FEATURE_THRESH_19_116": value  <= -0.00113433704245835543;
            "FEATURE_THRESH_19_117": value  <= 0.01681699976325039952;
            "FEATURE_THRESH_19_118": value  <= 0.00505351787433028221;
            "FEATURE_THRESH_19_119": value  <= -0.00458747101947665215;
            "FEATURE_THRESH_19_120": value  <= 0.00168824603315442801;
            "FEATURE_THRESH_19_121": value  <= -0.00165540003217756748;
            "FEATURE_THRESH_19_122": value  <= -0.01937380060553550026;
            "FEATURE_THRESH_19_123": value  <= 0.01037445012480020003;
            "FEATURE_THRESH_19_124": value  <= 0.00014973050565458834;
            "FEATURE_THRESH_19_125": value  <= -0.04298193007707599989;
            "FEATURE_THRESH_19_126": value  <= 0.00830659363418817520;
            "FEATURE_THRESH_19_127": value  <= -0.00412857905030250549;
            "FEATURE_THRESH_19_128": value  <= 0.00173994200304150581;
            "FEATURE_THRESH_19_129": value  <= 0.00011739750334527344;
            "FEATURE_THRESH_19_130": value  <= 0.00018585780344437808;
            "FEATURE_THRESH_19_131": value  <= 0.00555876921862363815;
            "FEATURE_THRESH_19_132": value  <= -0.00798515602946281433;
            "FEATURE_THRESH_19_133": value  <= 0.00060594122624024749;
            "FEATURE_THRESH_19_134": value  <= -0.00022983040253166109;
            "FEATURE_THRESH_19_135": value  <= 0.00043740210821852088;
            "FEATURE_THRESH_19_136": value  <= 0.00029482020181603730;
            "FEATURE_THRESH_19_137": value  <= 0.01031265966594220075;
            "FEATURE_THRESH_19_138": value  <= -0.00772411096841096878;
            "FEATURE_THRESH_19_139": value  <= -0.00467972084879875183;
            "FEATURE_THRESH_19_140": value  <= -0.00507554598152637482;
            "FEATURE_THRESH_19_141": value  <= 0.00224797404371201992;
            "FEATURE_THRESH_19_142": value  <= 0.00083327008178457618;
            "FEATURE_THRESH_19_143": value  <= -0.04127933084964750116;
            "FEATURE_THRESH_19_144": value  <= -0.00050930189900100231;
            "FEATURE_THRESH_19_145": value  <= 0.00125687802210450172;
            "FEATURE_THRESH_19_146": value  <= 0.00800484977662563324;
            "FEATURE_THRESH_19_147": value  <= -0.00118793000001460314;
            "FEATURE_THRESH_19_148": value  <= 0.00061948952497914433;
            "FEATURE_THRESH_19_149": value  <= 0.00668298592790961266;
            "FEATURE_THRESH_19_150": value  <= -0.00370623404160141945;
            "FEATURE_THRESH_19_151": value  <= -0.03973941132426259820;
            "FEATURE_THRESH_19_152": value  <= 0.00140850094612687826;
            "FEATURE_THRESH_19_153": value  <= 0.00039322688826359808;
            "FEATURE_THRESH_19_154": value  <= -0.00189798197243362665;
            "FEATURE_THRESH_19_155": value  <= -0.01397044025361540015;
            "FEATURE_THRESH_19_156": value  <= -0.10100819915533069959;
            "FEATURE_THRESH_19_157": value  <= -0.01734692044556139859;
            "FEATURE_THRESH_19_158": value  <= 0.00015619759506080300;
            "FEATURE_THRESH_19_159": value  <= 0.13438929617404940520;
            "FEATURE_THRESH_19_160": value  <= -0.02458224073052410127;
            "FEATURE_THRESH_19_161": value  <= -0.00385537208057940006;
            "FEATURE_THRESH_19_162": value  <= -0.00231652497313916683;
            "FEATURE_THRESH_19_163": value  <= -0.00485181203112006187;
            "FEATURE_THRESH_19_164": value  <= 0.00246999389491975307;
            "FEATURE_THRESH_19_165": value  <= 0.04549695923924450269;
            "FEATURE_THRESH_19_166": value  <= -0.02031959965825079831;
            "FEATURE_THRESH_19_167": value  <= 0.00026994998916052282;
            "FEATURE_THRESH_19_168": value  <= -0.00182326999492943287;
            "FEATURE_THRESH_19_169": value  <= -0.00630157906562089920;
            "FEATURE_THRESH_19_170": value  <= -0.00024139499873854220;
            "FEATURE_THRESH_19_171": value  <= -0.00103303696960210800;
            "FEATURE_THRESH_19_172": value  <= 0.00018041160365100950;
            "FEATURE_THRESH_19_173": value  <= -0.06140786036849019830;
            "FEATURE_THRESH_19_174": value  <= -0.06954391300678250398;
            "FEATURE_THRESH_19_175": value  <= -0.07054266333580019865;
            "FEATURE_THRESH_19_176": value  <= 0.00244237994775176048;
            "FEATURE_THRESH_19_177": value  <= 0.00154943496454507113;
            "FEATURE_THRESH_19_178": value  <= -0.02391421981155869916;
            "FEATURE_THRESH_19_179": value  <= -0.01245369017124180015;
            "FEATURE_THRESH_19_180": value  <= -0.00020760179904755205;
            "FEATURE_THRESH_19_181": value  <= 0.00002978108022944071;
            "FEATURE_THRESH_20_0": value  <= 0.01177274994552139978;
            "FEATURE_THRESH_20_1": value  <= 0.02703757025301459921;
            "FEATURE_THRESH_20_2": value  <= -0.00003641950024757534;
            "FEATURE_THRESH_20_3": value  <= 0.00199954095296561718;
            "FEATURE_THRESH_20_4": value  <= 0.00452783005312085152;
            "FEATURE_THRESH_20_5": value  <= 0.00047890920541249216;
            "FEATURE_THRESH_20_6": value  <= 0.00117209204472601414;
            "FEATURE_THRESH_20_7": value  <= 0.00095305702416226268;
            "FEATURE_THRESH_20_8": value  <= 0.00001509915000497131;
            "FEATURE_THRESH_20_9": value  <= -0.00060817901976406574;
            "FEATURE_THRESH_20_10": value  <= 0.00332245207391679287;
            "FEATURE_THRESH_20_11": value  <= -0.00110374903306365013;
            "FEATURE_THRESH_20_12": value  <= -0.00143502699211239815;
            "FEATURE_THRESH_20_13": value  <= 0.00207673991098999977;
            "FEATURE_THRESH_20_14": value  <= -0.00016412809782195836;
            "FEATURE_THRESH_20_15": value  <= 0.00883024372160434723;
            "FEATURE_THRESH_20_16": value  <= -0.01055207010358569925;
            "FEATURE_THRESH_20_17": value  <= -0.00227316003292798996;
            "FEATURE_THRESH_20_18": value  <= -0.00084786332445219159;
            "FEATURE_THRESH_20_19": value  <= 0.00120813597459346056;
            "FEATURE_THRESH_20_20": value  <= 0.00265127304010093212;
            "FEATURE_THRESH_20_21": value  <= -0.00110124796628952026;
            "FEATURE_THRESH_20_22": value  <= 0.00049561518244445324;
            "FEATURE_THRESH_20_23": value  <= -0.04390177130699159797;
            "FEATURE_THRESH_20_24": value  <= 0.03469035029411320081;
            "FEATURE_THRESH_20_25": value  <= -0.00274421903304755688;
            "FEATURE_THRESH_20_26": value  <= 0.00333165889605879784;
            "FEATURE_THRESH_20_27": value  <= -0.02004457078874110135;
            "FEATURE_THRESH_20_28": value  <= 0.00134920305572450161;
            "FEATURE_THRESH_20_29": value  <= 0.00297020189464092255;
            "FEATURE_THRESH_20_30": value  <= 0.00630399817600846291;
            "FEATURE_THRESH_20_31": value  <= -0.01293659023940560079;
            "FEATURE_THRESH_20_32": value  <= 0.00401487294584512711;
            "FEATURE_THRESH_20_33": value  <= -0.00264016794972121716;
            "FEATURE_THRESH_20_34": value  <= 0.01391843985766169980;
            "FEATURE_THRESH_20_35": value  <= -0.00045087869511917233;
            "FEATURE_THRESH_20_36": value  <= 0.00025384349282830954;
            "FEATURE_THRESH_20_37": value  <= 0.00227100006304681301;
            "FEATURE_THRESH_20_38": value  <= 0.00241207797080278397;
            "FEATURE_THRESH_20_39": value  <= -0.00003602567085181363;
            "FEATURE_THRESH_20_40": value  <= -0.00749055296182632446;
            "FEATURE_THRESH_20_41": value  <= -0.01751312054693699924;
            "FEATURE_THRESH_20_42": value  <= 0.14281630516052248869;
            "FEATURE_THRESH_20_43": value  <= 0.00553452689200639725;
            "FEATURE_THRESH_20_44": value  <= -0.00096323591424152255;
            "FEATURE_THRESH_20_45": value  <= -0.00203700107522308826;
            "FEATURE_THRESH_20_46": value  <= 0.00166148296557366848;
            "FEATURE_THRESH_20_47": value  <= -0.00311880907975137234;
            "FEATURE_THRESH_20_48": value  <= -0.00640006177127361298;
            "FEATURE_THRESH_20_49": value  <= 0.00031319601112045348;
            "FEATURE_THRESH_20_50": value  <= -0.01822209917008879923;
            "FEATURE_THRESH_20_51": value  <= 0.00879692472517490387;
            "FEATURE_THRESH_20_52": value  <= -0.00423950701951980591;
            "FEATURE_THRESH_20_53": value  <= 0.00970862712711095810;
            "FEATURE_THRESH_20_54": value  <= -0.00399341713637113571;
            "FEATURE_THRESH_20_55": value  <= -0.01678505912423130034;
            "FEATURE_THRESH_20_56": value  <= 0.01827209070324899848;
            "FEATURE_THRESH_20_57": value  <= 0.00568728381767868996;
            "FEATURE_THRESH_20_58": value  <= -0.00107390398625284433;
            "FEATURE_THRESH_20_59": value  <= -0.00370938703417778015;
            "FEATURE_THRESH_20_60": value  <= -0.00021110709349159151;
            "FEATURE_THRESH_20_61": value  <= 0.00106701394543051720;
            "FEATURE_THRESH_20_62": value  <= 0.00359430210664868355;
            "FEATURE_THRESH_20_63": value  <= -0.00517760310322046280;
            "FEATURE_THRESH_20_64": value  <= -0.00025414369883947074;
            "FEATURE_THRESH_20_65": value  <= 0.00635225605219602585;
            "FEATURE_THRESH_20_66": value  <= -0.00044205080484971404;
            "FEATURE_THRESH_20_67": value  <= 0.00074488727841526270;
            "FEATURE_THRESH_20_68": value  <= -0.00351163791492581367;
            "FEATURE_THRESH_20_69": value  <= -0.01254091039299960048;
            "FEATURE_THRESH_20_70": value  <= 0.00949318520724773407;
            "FEATURE_THRESH_20_71": value  <= 0.01296115014702079946;
            "FEATURE_THRESH_20_72": value  <= 0.00472094491124153137;
            "FEATURE_THRESH_20_73": value  <= -0.00231190794147551060;
            "FEATURE_THRESH_20_74": value  <= -0.00282622990198433399;
            "FEATURE_THRESH_20_75": value  <= -0.00143113394733518362;
            "FEATURE_THRESH_20_76": value  <= 0.00193783105351030827;
            "FEATURE_THRESH_20_77": value  <= 0.00026343559147790074;
            "FEATURE_THRESH_20_78": value  <= 0.00078257522545754910;
            "FEATURE_THRESH_20_79": value  <= -0.01955044083297249879;
            "FEATURE_THRESH_20_80": value  <= 0.00043914958951063454;
            "FEATURE_THRESH_20_81": value  <= 0.02145200036466119939;
            "FEATURE_THRESH_20_82": value  <= 0.00058973580598831177;
            "FEATURE_THRESH_20_83": value  <= -0.02615761011838909841;
            "FEATURE_THRESH_20_84": value  <= -0.01395986042916770066;
            "FEATURE_THRESH_20_85": value  <= -0.00636990182101726532;
            "FEATURE_THRESH_20_86": value  <= -0.00856138207018375397;
            "FEATURE_THRESH_20_87": value  <= 0.00096622901037335396;
            "FEATURE_THRESH_20_88": value  <= 0.00076550268568098545;
            "FEATURE_THRESH_20_89": value  <= -0.00818333402276039124;
            "FEATURE_THRESH_20_90": value  <= -0.00939769390970468521;
            "FEATURE_THRESH_20_91": value  <= 0.00480289803817868233;
            "FEATURE_THRESH_20_92": value  <= -0.00356805697083473206;
            "FEATURE_THRESH_20_93": value  <= 0.00407331204041838646;
            "FEATURE_THRESH_20_94": value  <= 0.00125681294593960047;
            "FEATURE_THRESH_20_95": value  <= -0.00290650106035172939;
            "FEATURE_THRESH_20_96": value  <= -0.00244093406945466995;
            "FEATURE_THRESH_20_97": value  <= 0.02483070082962509847;
            "FEATURE_THRESH_20_98": value  <= -0.04885400831699369950;
            "FEATURE_THRESH_20_99": value  <= -0.00161103799473494291;
            "FEATURE_THRESH_20_100": value  <= -0.09700947999954219469;
            "FEATURE_THRESH_20_101": value  <= 0.00112092401832342148;
            "FEATURE_THRESH_20_102": value  <= -0.00130640901625156403;
            "FEATURE_THRESH_20_103": value  <= 0.00045771620352752507;
            "FEATURE_THRESH_20_104": value  <= -0.00063149951165542006;
            "FEATURE_THRESH_20_105": value  <= 0.00014505970466416329;
            "FEATURE_THRESH_20_106": value  <= -0.01647455058991910068;
            "FEATURE_THRESH_20_107": value  <= 0.01336957979947329955;
            "FEATURE_THRESH_20_108": value  <= 0.00010271780047332868;
            "FEATURE_THRESH_20_109": value  <= -0.00553115596994757652;
            "FEATURE_THRESH_20_110": value  <= -0.00261870492249727249;
            "FEATURE_THRESH_20_111": value  <= 0.00508342683315277100;
            "FEATURE_THRESH_20_112": value  <= 0.07981815934181210603;
            "FEATURE_THRESH_20_113": value  <= -0.09922658652067180285;
            "FEATURE_THRESH_20_114": value  <= -0.00065174017800018191;
            "FEATURE_THRESH_20_115": value  <= -0.01899684965610499987;
            "FEATURE_THRESH_20_116": value  <= 0.01734689995646479868;
            "FEATURE_THRESH_20_117": value  <= 0.00055082101607695222;
            "FEATURE_THRESH_20_118": value  <= 0.00200560502707958221;
            "FEATURE_THRESH_20_119": value  <= -0.00776881910860538483;
            "FEATURE_THRESH_20_120": value  <= 0.05087827891111369738;
            "FEATURE_THRESH_20_121": value  <= -0.00229017809033393860;
            "FEATURE_THRESH_20_122": value  <= -0.00015715380141045898;
            "FEATURE_THRESH_20_123": value  <= 0.10519240051507949829;
            "FEATURE_THRESH_20_124": value  <= 0.00271989195607602596;
            "FEATURE_THRESH_20_125": value  <= 0.04833777993917470067;
            "FEATURE_THRESH_20_126": value  <= 0.00095703761326149106;
            "FEATURE_THRESH_20_127": value  <= -0.02537125907838340064;
            "FEATURE_THRESH_20_128": value  <= 0.05245795100927350130;
            "FEATURE_THRESH_20_129": value  <= -0.01236562989652159952;
            "FEATURE_THRESH_20_130": value  <= -0.14589719474315640535;
            "FEATURE_THRESH_20_131": value  <= -0.01590860076248649946;
            "FEATURE_THRESH_20_132": value  <= 0.00039486068999394774;
            "FEATURE_THRESH_20_133": value  <= -0.00524540012702345848;
            "FEATURE_THRESH_20_134": value  <= -0.00504217995330691338;
            "FEATURE_THRESH_20_135": value  <= 0.00298121897503733635;
            "FEATURE_THRESH_20_136": value  <= -0.00728843081742525101;
            "FEATURE_THRESH_20_137": value  <= 0.00150943500921130180;
            "FEATURE_THRESH_20_138": value  <= -0.00933407992124557495;
            "FEATURE_THRESH_20_139": value  <= 0.02866714075207709919;
            "FEATURE_THRESH_20_140": value  <= 0.17019680142402648926;
            "FEATURE_THRESH_20_141": value  <= -0.00326144788414239883;
            "FEATURE_THRESH_20_142": value  <= 0.00055769277969375253;
            "FEATURE_THRESH_20_143": value  <= 0.36258339881896972656;
            "FEATURE_THRESH_20_144": value  <= -0.01161513011902570031;
            "FEATURE_THRESH_20_145": value  <= -0.00407951977103948593;
            "FEATURE_THRESH_20_146": value  <= 0.00057204300537705421;
            "FEATURE_THRESH_20_147": value  <= 0.00067543348995968699;
            "FEATURE_THRESH_20_148": value  <= 0.00063295697327703238;
            "FEATURE_THRESH_20_149": value  <= 0.00124353205319494009;
            "FEATURE_THRESH_20_150": value  <= -0.00473638577386736870;
            "FEATURE_THRESH_20_151": value  <= -0.00646584620699286461;
            "FEATURE_THRESH_20_152": value  <= 0.00035017321351915598;
            "FEATURE_THRESH_20_153": value  <= 0.00015754920605104417;
            "FEATURE_THRESH_20_154": value  <= 0.00997743662446737289;
            "FEATURE_THRESH_20_155": value  <= -0.00041464529931545258;
            "FEATURE_THRESH_20_156": value  <= -0.00035888899583369493;
            "FEATURE_THRESH_20_157": value  <= 0.00040463250479660928;
            "FEATURE_THRESH_20_158": value  <= -0.00082184787606820464;
            "FEATURE_THRESH_20_159": value  <= 0.00594674190506339073;
            "FEATURE_THRESH_20_160": value  <= -0.02175338938832279898;
            "FEATURE_THRESH_20_161": value  <= -0.01454037986695769918;
            "FEATURE_THRESH_20_162": value  <= -0.04051076993346210131;
            "FEATURE_THRESH_20_163": value  <= -0.00058458268176764250;
            "FEATURE_THRESH_20_164": value  <= 0.00551518006250262260;
            "FEATURE_THRESH_20_165": value  <= -0.00606262218207120895;
            "FEATURE_THRESH_20_166": value  <= 0.09453584253787990221;
            "FEATURE_THRESH_20_167": value  <= 0.00473150517791509628;
            "FEATURE_THRESH_20_168": value  <= -0.00052571471314877272;
            "FEATURE_THRESH_20_169": value  <= -0.00254640495404601097;
            "FEATURE_THRESH_20_170": value  <= -0.02607568912208079945;
            "FEATURE_THRESH_20_171": value  <= -0.00547797093167901039;
            "FEATURE_THRESH_20_172": value  <= 0.00513377413153648376;
            "FEATURE_THRESH_20_173": value  <= 0.00047944980906322598;
            "FEATURE_THRESH_20_174": value  <= -0.00211140792816877365;
            "FEATURE_THRESH_20_175": value  <= -0.01317999046295880057;
            "FEATURE_THRESH_20_176": value  <= -0.00479680998250842094;
            "FEATURE_THRESH_20_177": value  <= 0.00674831680953502655;
            "FEATURE_THRESH_20_178": value  <= 0.00146233697887510061;
            "FEATURE_THRESH_20_179": value  <= 0.00476451590657234192;
            "FEATURE_THRESH_20_180": value  <= 0.00680666603147983551;
            "FEATURE_THRESH_20_181": value  <= 0.00366086210124194622;
            "FEATURE_THRESH_20_182": value  <= 0.02144964039325709948;
            "FEATURE_THRESH_20_183": value  <= 0.00416789017617702484;
            "FEATURE_THRESH_20_184": value  <= 0.00864675641059875488;
            "FEATURE_THRESH_20_185": value  <= -0.00036114078829996288;
            "FEATURE_THRESH_20_186": value  <= 0.00108087295666337013;
            "FEATURE_THRESH_20_187": value  <= 0.00577199598774313927;
            "FEATURE_THRESH_20_188": value  <= 0.00157207704614847898;
            "FEATURE_THRESH_20_189": value  <= -0.00193078594747930765;
            "FEATURE_THRESH_20_190": value  <= -0.00789262726902961731;
            "FEATURE_THRESH_20_191": value  <= -0.00222246791236102581;
            "FEATURE_THRESH_20_192": value  <= 0.00190119899343699217;
            "FEATURE_THRESH_20_193": value  <= 0.00275761191733181477;
            "FEATURE_THRESH_20_194": value  <= 0.00517874490469694138;
            "FEATURE_THRESH_20_195": value  <= -0.00090273341629654169;
            "FEATURE_THRESH_20_196": value  <= 0.00517979590222239494;
            "FEATURE_THRESH_20_197": value  <= -0.01011400017887350081;
            "FEATURE_THRESH_20_198": value  <= -0.01861706003546709925;
            "FEATURE_THRESH_20_199": value  <= 0.00592259597033262253;
            "FEATURE_THRESH_20_200": value  <= -0.00629450799897313118;
            "FEATURE_THRESH_20_201": value  <= 0.00653530191630125046;
            "FEATURE_THRESH_20_202": value  <= 0.00108783994801342487;
            "FEATURE_THRESH_20_203": value  <= -0.02254224009811879939;
            "FEATURE_THRESH_20_204": value  <= -0.00300656608305871487;
            "FEATURE_THRESH_20_205": value  <= 0.00747412722557783127;
            "FEATURE_THRESH_20_206": value  <= 0.02616232074797150003;
            "FEATURE_THRESH_20_207": value  <= 0.00094352738233283162;
            "FEATURE_THRESH_20_208": value  <= 0.03336324170231819847;
            "FEATURE_THRESH_20_209": value  <= -0.01511865016072990071;
            "FEATURE_THRESH_20_210": value  <= 0.00098648946732282639;
            "FEATURE_THRESH_21_0": value  <= -0.09515079855918880114;
            "FEATURE_THRESH_21_1": value  <= 0.00627023400738835335;
            "FEATURE_THRESH_21_2": value  <= 0.00030018089455552399;
            "FEATURE_THRESH_21_3": value  <= 0.00117574096657335758;
            "FEATURE_THRESH_21_4": value  <= 0.00004423526843311266;
            "FEATURE_THRESH_21_5": value  <= -0.00002993692032760010;
            "FEATURE_THRESH_21_6": value  <= 0.00300731998868286610;
            "FEATURE_THRESH_21_7": value  <= -0.01051388960331679952;
            "FEATURE_THRESH_21_8": value  <= 0.00834768265485763550;
            "FEATURE_THRESH_21_9": value  <= -0.00314922700636088848;
            "FEATURE_THRESH_21_10": value  <= -0.00001443564997316571;
            "FEATURE_THRESH_21_11": value  <= -0.00042855090578086674;
            "FEATURE_THRESH_21_12": value  <= 0.00015062429883982986;
            "FEATURE_THRESH_21_13": value  <= 0.07155983150005340576;
            "FEATURE_THRESH_21_14": value  <= 0.00084095180500298738;
            "FEATURE_THRESH_21_15": value  <= 0.06298650056123729357;
            "FEATURE_THRESH_21_16": value  <= -0.00337986298836767673;
            "FEATURE_THRESH_21_17": value  <= -0.00011810739670181647;
            "FEATURE_THRESH_21_18": value  <= -0.00054505601292476058;
            "FEATURE_THRESH_21_19": value  <= -0.00184549100231379271;
            "FEATURE_THRESH_21_20": value  <= -0.00043832371011376381;
            "FEATURE_THRESH_21_21": value  <= -0.00240008300170302391;
            "FEATURE_THRESH_21_22": value  <= -0.09879574179649350252;
            "FEATURE_THRESH_21_23": value  <= 0.00317982397973537445;
            "FEATURE_THRESH_21_24": value  <= 0.00032406419632025063;
            "FEATURE_THRESH_21_25": value  <= -0.03254725039005280235;
            "FEATURE_THRESH_21_26": value  <= -0.00775611307471990585;
            "FEATURE_THRESH_21_27": value  <= 0.01602724939584729974;
            "FEATURE_THRESH_21_28": value  <= 0.00000710023505234858;
            "FEATURE_THRESH_21_29": value  <= 0.00734228082001209259;
            "FEATURE_THRESH_21_30": value  <= -0.00169702805578708649;
            "FEATURE_THRESH_21_31": value  <= 0.00241182604804635048;
            "FEATURE_THRESH_21_32": value  <= -0.00553009379655122757;
            "FEATURE_THRESH_21_33": value  <= -0.00264787301421165466;
            "FEATURE_THRESH_21_34": value  <= 0.01129562966525549973;
            "FEATURE_THRESH_21_35": value  <= -0.00066952878842130303;
            "FEATURE_THRESH_21_36": value  <= 0.00144106801599264145;
            "FEATURE_THRESH_21_37": value  <= 0.00246378709562122822;
            "FEATURE_THRESH_21_38": value  <= 0.00033114518737420440;
            "FEATURE_THRESH_21_39": value  <= -0.03355726972222330268;
            "FEATURE_THRESH_21_40": value  <= 0.01853941939771179895;
            "FEATURE_THRESH_21_41": value  <= -0.00029698139405809343;
            "FEATURE_THRESH_21_42": value  <= -0.00045577259152196348;
            "FEATURE_THRESH_21_43": value  <= -0.01015898026525969937;
            "FEATURE_THRESH_21_44": value  <= -0.00002241382935608272;
            "FEATURE_THRESH_21_45": value  <= 0.00007203496352303773;
            "FEATURE_THRESH_21_46": value  <= -0.00692672096192836761;
            "FEATURE_THRESH_21_47": value  <= -0.00769978389143943787;
            "FEATURE_THRESH_21_48": value  <= -0.00731305498629808426;
            "FEATURE_THRESH_21_49": value  <= 0.00196505896747112274;
            "FEATURE_THRESH_21_50": value  <= 0.00716476002708077431;
            "FEATURE_THRESH_21_51": value  <= -0.02407863922417160032;
            "FEATURE_THRESH_21_52": value  <= -0.02102796919643879978;
            "FEATURE_THRESH_21_53": value  <= 0.00036017020465806127;
            "FEATURE_THRESH_21_54": value  <= -0.01721972972154620085;
            "FEATURE_THRESH_21_55": value  <= -0.00786721426993608475;
            "FEATURE_THRESH_21_56": value  <= -0.00044777389848604798;
            "FEATURE_THRESH_21_57": value  <= 0.00554860103875398636;
            "FEATURE_THRESH_21_58": value  <= -0.00694611482322216034;
            "FEATURE_THRESH_21_59": value  <= 0.00013569870498031378;
            "FEATURE_THRESH_21_60": value  <= -0.04588025063276290200;
            "FEATURE_THRESH_21_61": value  <= -0.02158256061375140103;
            "FEATURE_THRESH_21_62": value  <= -0.02020953968167309850;
            "FEATURE_THRESH_21_63": value  <= 0.00584967108443379402;
            "FEATURE_THRESH_21_64": value  <= -0.00005747637987951749;
            "FEATURE_THRESH_21_65": value  <= -0.00115131004713475704;
            "FEATURE_THRESH_21_66": value  <= 0.00198628311045467854;
            "FEATURE_THRESH_21_67": value  <= -0.00527195120230317116;
            "FEATURE_THRESH_21_68": value  <= 0.00126626994460821152;
            "FEATURE_THRESH_21_69": value  <= -0.00629194406792521477;
            "FEATURE_THRESH_21_70": value  <= 0.00067360111279413104;
            "FEATURE_THRESH_21_71": value  <= -0.00105234503280371428;
            "FEATURE_THRESH_21_72": value  <= -0.00044216238893568516;
            "FEATURE_THRESH_21_73": value  <= 0.00117479404434561729;
            "FEATURE_THRESH_21_74": value  <= 0.00524574378505349159;
            "FEATURE_THRESH_21_75": value  <= -0.02453972026705740148;
            "FEATURE_THRESH_21_76": value  <= 0.00073793041519820690;
            "FEATURE_THRESH_21_77": value  <= 0.00142337998840957880;
            "FEATURE_THRESH_21_78": value  <= -0.00241491105407476425;
            "FEATURE_THRESH_21_79": value  <= -0.00121652998495846987;
            "FEATURE_THRESH_21_80": value  <= -0.00124388094991445541;
            "FEATURE_THRESH_21_81": value  <= 0.00619427394121885300;
            "FEATURE_THRESH_21_82": value  <= -0.00166071695275604725;
            "FEATURE_THRESH_21_83": value  <= -0.02731625922024250031;
            "FEATURE_THRESH_21_84": value  <= -0.00158455700147897005;
            "FEATURE_THRESH_21_85": value  <= -0.00155147397890686989;
            "FEATURE_THRESH_21_86": value  <= 0.00038446558755822480;
            "FEATURE_THRESH_21_87": value  <= -0.01467225980013609973;
            "FEATURE_THRESH_21_88": value  <= 0.00816088821738958359;
            "FEATURE_THRESH_21_89": value  <= 0.00111216597724705935;
            "FEATURE_THRESH_21_90": value  <= -0.00726037705317139626;
            "FEATURE_THRESH_21_91": value  <= -0.00024046430189628154;
            "FEATURE_THRESH_21_92": value  <= -0.00023348190006799996;
            "FEATURE_THRESH_21_93": value  <= 0.00557364802807569504;
            "FEATURE_THRESH_21_94": value  <= 0.03062376938760279915;
            "FEATURE_THRESH_21_95": value  <= 0.00092074798885732889;
            "FEATURE_THRESH_21_96": value  <= -0.00004355073906481267;
            "FEATURE_THRESH_21_97": value  <= -0.00664527108892798424;
            "FEATURE_THRESH_21_98": value  <= 0.04322199895977969775;
            "FEATURE_THRESH_21_99": value  <= 0.00223317695781588554;
            "FEATURE_THRESH_21_100": value  <= 0.00318297394551336765;
            "FEATURE_THRESH_21_101": value  <= -0.00018027749320026487;
            "FEATURE_THRESH_21_102": value  <= -0.00529346894472837448;
            "FEATURE_THRESH_21_103": value  <= 0.00127509597223252058;
            "FEATURE_THRESH_21_104": value  <= 0.00433853222057223320;
            "FEATURE_THRESH_21_105": value  <= 0.00852507445961236954;
            "FEATURE_THRESH_21_106": value  <= -0.00094266352243721485;
            "FEATURE_THRESH_21_107": value  <= 0.00136096600908786058;
            "FEATURE_THRESH_21_108": value  <= 0.00044782509212382138;
            "FEATURE_THRESH_21_109": value  <= 0.00133600505068898201;
            "FEATURE_THRESH_21_110": value  <= -0.00060967548051849008;
            "FEATURE_THRESH_21_111": value  <= -0.00236567808315157890;
            "FEATURE_THRESH_21_112": value  <= 0.00107343401759862900;
            "FEATURE_THRESH_21_113": value  <= 0.00219233590178191662;
            "FEATURE_THRESH_21_114": value  <= 0.00549686187878251076;
            "FEATURE_THRESH_21_115": value  <= -0.07536882162094120374;
            "FEATURE_THRESH_21_116": value  <= 0.02513447031378749849;
            "FEATURE_THRESH_21_117": value  <= -0.00002935859993158374;
            "FEATURE_THRESH_21_118": value  <= -0.00058355910005047917;
            "FEATURE_THRESH_21_119": value  <= -0.00266394508071243763;
            "FEATURE_THRESH_21_120": value  <= -0.00138040899764746428;
            "FEATURE_THRESH_21_121": value  <= 0.00123132194858044386;
            "FEATURE_THRESH_21_122": value  <= -0.00001464417982788291;
            "FEATURE_THRESH_21_123": value  <= -0.01281880959868430050;
            "FEATURE_THRESH_21_124": value  <= 0.02285218983888629915;
            "FEATURE_THRESH_21_125": value  <= 0.00082305970136076212;
            "FEATURE_THRESH_21_126": value  <= 0.01277012005448339982;
            "FEATURE_THRESH_21_127": value  <= -0.05005151033401489952;
            "FEATURE_THRESH_21_128": value  <= 0.01577527076005939832;
            "FEATURE_THRESH_21_129": value  <= -0.01850162073969839963;
            "FEATURE_THRESH_21_130": value  <= 0.00246262503787875175;
            "FEATURE_THRESH_21_131": value  <= 0.06291616708040240202;
            "FEATURE_THRESH_21_132": value  <= -0.00002164850047847722;
            "FEATURE_THRESH_21_133": value  <= 0.00211809901520609856;
            "FEATURE_THRESH_21_134": value  <= -0.01663489080965519992;
            "FEATURE_THRESH_21_135": value  <= -0.00288994703441858292;
            "FEATURE_THRESH_21_136": value  <= 0.07678326219320300017;
            "FEATURE_THRESH_21_137": value  <= 0.00391706777736544609;
            "FEATURE_THRESH_21_138": value  <= -0.07267060130834579468;
            "FEATURE_THRESH_21_139": value  <= 0.54039502143859863281;
            "FEATURE_THRESH_21_140": value  <= 0.00295100198127329350;
            "FEATURE_THRESH_21_141": value  <= 0.00345083698630332947;
            "FEATURE_THRESH_21_142": value  <= -0.00042077939724549651;
            "FEATURE_THRESH_21_143": value  <= 0.00330510502681136131;
            "FEATURE_THRESH_21_144": value  <= 0.00047735060798004270;
            "FEATURE_THRESH_21_145": value  <= -0.02592851035296920084;
            "FEATURE_THRESH_21_146": value  <= -0.00297297909855842590;
            "FEATURE_THRESH_21_147": value  <= 0.00585083290934562683;
            "FEATURE_THRESH_21_148": value  <= -0.04596751928329469855;
            "FEATURE_THRESH_21_149": value  <= 0.15585960447788241301;
            "FEATURE_THRESH_21_150": value  <= 0.01516482979059220054;
            "FEATURE_THRESH_21_151": value  <= -0.00106042495463043451;
            "FEATURE_THRESH_21_152": value  <= 0.00664762919768691063;
            "FEATURE_THRESH_21_153": value  <= -0.01223113015294080043;
            "FEATURE_THRESH_21_154": value  <= 0.00565288821235299110;
            "FEATURE_THRESH_21_155": value  <= 0.00129778299015015364;
            "FEATURE_THRESH_21_156": value  <= 0.01078158989548680044;
            "FEATURE_THRESH_21_157": value  <= 0.00286547793075442314;
            "FEATURE_THRESH_21_158": value  <= 0.00286634289659559727;
            "FEATURE_THRESH_21_159": value  <= -0.00519833201542496681;
            "FEATURE_THRESH_21_160": value  <= 0.00537399901077151299;
            "FEATURE_THRESH_21_161": value  <= -0.01464152988046409955;
            "FEATURE_THRESH_21_162": value  <= -0.00001504258034401573;
            "FEATURE_THRESH_21_163": value  <= -0.00011875660129589960;
            "FEATURE_THRESH_21_164": value  <= 0.01699553057551380156;
            "FEATURE_THRESH_21_165": value  <= -0.03509594127535820007;
            "FEATURE_THRESH_21_166": value  <= 0.00242173508740961552;
            "FEATURE_THRESH_21_167": value  <= -0.00096340337768197060;
            "FEATURE_THRESH_21_168": value  <= 0.00016391130338888615;
            "FEATURE_THRESH_21_169": value  <= -0.02114146016538140035;
            "FEATURE_THRESH_21_170": value  <= 0.00087775202700868249;
            "FEATURE_THRESH_21_171": value  <= -0.02794392034411430012;
            "FEATURE_THRESH_21_172": value  <= 0.00672973785549402237;
            "FEATURE_THRESH_21_173": value  <= 0.02328103967010970027;
            "FEATURE_THRESH_21_174": value  <= -0.01164497993886469927;
            "FEATURE_THRESH_21_175": value  <= 0.01576430909335610128;
            "FEATURE_THRESH_21_176": value  <= -0.00136114796623587608;
            "FEATURE_THRESH_21_177": value  <= -0.00081522337859496474;
            "FEATURE_THRESH_21_178": value  <= -0.00060066272271797061;
            "FEATURE_THRESH_21_179": value  <= 0.00049715518252924085;
            "FEATURE_THRESH_21_180": value  <= 0.00234753708355128765;
            "FEATURE_THRESH_21_181": value  <= -0.00892615690827369690;
            "FEATURE_THRESH_21_182": value  <= -0.01391991041600700030;
            "FEATURE_THRESH_21_183": value  <= 0.00102099496871232986;
            "FEATURE_THRESH_21_184": value  <= -0.00274416292086243629;
            "FEATURE_THRESH_21_185": value  <= -0.01620013080537319877;
            "FEATURE_THRESH_21_186": value  <= 0.00433319807052612305;
            "FEATURE_THRESH_21_187": value  <= 0.00058497930876910686;
            "FEATURE_THRESH_21_188": value  <= -0.00224664504639804363;
            "FEATURE_THRESH_21_189": value  <= 0.00231460994109511375;
            "FEATURE_THRESH_21_190": value  <= 0.00876791216433048248;
            "FEATURE_THRESH_21_191": value  <= -0.00022448020172305405;
            "FEATURE_THRESH_21_192": value  <= -0.00743360212072730064;
            "FEATURE_THRESH_21_193": value  <= -0.00231892406009137630;
            "FEATURE_THRESH_21_194": value  <= -0.00210421788506209850;
            "FEATURE_THRESH_21_195": value  <= 0.00046034841216169298;
            "FEATURE_THRESH_21_196": value  <= 0.00105476297903805971;
            "FEATURE_THRESH_21_197": value  <= 0.00087148818420246243;
            "FEATURE_THRESH_21_198": value  <= 0.00033364820410497487;
            "FEATURE_THRESH_21_199": value  <= -0.00148532504681497812;
            "FEATURE_THRESH_21_200": value  <= 0.00302516203373670578;
            "FEATURE_THRESH_21_201": value  <= 0.00502807414159178734;
            "FEATURE_THRESH_21_202": value  <= -0.00058164511574432254;
            "FEATURE_THRESH_21_203": value  <= 0.04514152929186820290;
            "FEATURE_THRESH_21_204": value  <= -0.00107956200372427702;
            "FEATURE_THRESH_21_205": value  <= 0.00015995999274309725;
            "FEATURE_THRESH_21_206": value  <= -0.01935927011072640161;
            "FEATURE_THRESH_21_207": value  <= 0.20725509524345400725;
            "FEATURE_THRESH_21_208": value  <= -0.00041953290929086506;
            "FEATURE_THRESH_21_209": value  <= 0.00225820695050060749;
            "FEATURE_THRESH_21_210": value  <= -0.00678112078458070755;
            "FEATURE_THRESH_21_211": value  <= 0.01115430984646080016;
            "FEATURE_THRESH_21_212": value  <= 0.04316243156790729868;

            default: value <= 0;

        endcase

    end

endmodule 
